PK   +��Xv_��9  	    cirkitFile.json�}�n$����?Q��gD�s��X;cc<�Y�����[��R�J嶷�ڗ�g��L�������mՎ��S]�<q���7~�z����6��C��9=|����zG����a����V__}���<�o���}�������z�뇤��ԍ�=��LnңwA�X�t�����5�ѭ��h6z���}�����Ao��C-�ޘj�zc�9�"荫�P��7��C-�ބj�z�9�"�MS͡Ao�j��Q�BY�, RY��T/��̢^.�!�E�`VC0�z��B� �?~��Kw���141(�Qn���OFY�L�1q�����[�,�%��Yԋn5����-��}���)S���̢^��!�`�[�٦^�����X�S�z_�,����Y�kv5ĶJ�Y�k����j�m7\͢~�l�u��Y��n5����jf�Z�+�z�`���?���ݾ/�|��=�>�Uݥ?Uu(tLgmf*�3[���̢^ë!�E��WC0�z���W���̢^ë!�E��WC0�z��`�	�zw���jfQ���̢^;�!�E�vVC0�z��_���̢^;����ʱ����jfQ���̢^w���M_[��e�z����]�,�5{�����Y���̢^�!�&��}5����jfQ��3��!�~��?�����!�Z�<�Q;��X�Fs���v���p�dw Wώ��ˎ�k;���a�q���bmeGXv�am簶��#,;�`m籶��#,;�`m����#,;��X�E����No������NoZ��Z����.�N��cw�#0���l?tt�/���GX~��2���2���/���i`��_�?�8���#0��{l?pā�G`~y�=�~�ˏ�����������`���,?��'-����ˏ�����������m�`��W8�K��À��?���/ou�`��_�\�8���#0���l?p���G`~��~��ˏ����7��������s{`���,?��'��4�����峒`���,?�o���w�,8j������Q���V�nu����o�jkq���
��jC�9c�Yp0��G`~��!��;/h�:�]i.p,7�y���r�a��_>K�8���#0�|
l?p,��G`~��>�~�Xˏ��r���8���#0��3l?p,��G`~9��~�$,?��y*���%a��_ΰ�����8|q��Łג���/g5�`��_���8���#0��Il?p���G`~9�~��ˏ��r���<8���#0��w�dּ1�֓r1X[���_��8��݆*g��,4x5S9�8�
Rk�ǃ�,?��Y���G=X~��[���i�ɴʛ�W.p+�t�(ӏ�\?Qȯ��QYV�"*u�~t�*8<H��������c-��<8���#0��G�D5t�"�^+;�I9���w�Ʃ�d�D��k�pT�U����Up�7�i��Gx�a��_�z�8���#0����D5bg�sug��\��!F����4%=U��T�U��J�j̭�Ã�x]+�׵���/gf��a��~+7���\�箮�qB̕ŏ��޻X���(���r��we��Ľ+�'�]Y���$m�َSܮ�^]3s�k���V�����R����yt�Վ���-_��fob\�E'9����r9�R��|e㛽�pm�ھ���G5�_jEE�tU6�������ǻ�Ǉ��Ǫ���Ǜ��4������m�����{k�/kNa�Ws�e�����G��G��N�8���b�T����y�:*Ǔ�T�ކ��E�^� g�qF\�Ϣ@fYZ��/+KQ�e;Fa�Ԙ�6?^���R����E��T
c��^��
��TZ�`V��8���TPY�j**��6y�)��3=�\�b_�����D!���p����v2�*
�S��=�[MS�al�b�]�z��E�����p��\�:K�E�O�x������~sѓ���0�#{;��)�P���-)jFK��x��.*~& ��Q5cb�n,D��j�z���ug�^T|��cC�o���/���Ρw�SSc8Ԛ��M{��Eŗ�>hc��
r�n0�W��H��0���Ӌ�����n�ڨF�]���Qm��fl�زC��,_R���ˀ�AQj�1�ߛ�YŰ}��7�Н�|I���a���<������6�o[�N��=�����;��0i�zC���6�K)�G��5��?��E��x�dm�'X3p�q��8�Siơo�y��ו_~z0��q�Zρ����fP��� �Y����ӹ���u*�M��̤��X7c�m�.�tN�J�/?]����e�g�h�W�����ɞ�|Q�sj��G7�������u���7f0�����zS�)x����&�쾭��kzbe�1�꽤��9���ʴL�K���k��R�l�sO/*~�G�����.�O�R=��!�vbύ�\{/*����Oڲ>8��&ͽt��0t���<������W\O��r�"�kת!�oH��4�����gZ\��NF��c������wj�c��O�kq%ŷO�۶���~3ܿ��z����m�������~\�~�m�F ���h;-�a�Na����FF ��n#�v�	�h�g���˂a�m�I$N�q��m�	7
i�I�	��o�nG��i����L�QH��K N0'����v��@�ڝ?�c����(���-'��7 �鸁�����Ws��8
i���	670G!��8�t��t��ۨ��[����v;�@�`:na:�B��a�`�q�q�62#Q���W�	6�0G!��0N0�0G!�$�0N0w0G!�d�0N0w0G!夝0N�9qܤ8L�l<�B�	a�`:�`:�Bʉa�`:�`:�B�	�`K?0�0F�&�`:�B�i�`�`:�a:�C���8Z��[ބ鸇�8
)$�q�"��G=Vr��8
)��q��x��8
)'q�q���LǗ���8��s���-u�a�Ԍ���-s���\v=��G�q%�$�Uo�s�Q�v��J"\��8,hW	�$�.�gk�X@�+�p�q��]���b, ��D��EĮ��]1��J"\��8�*hW	�$�Uo�3��Q�v��J"\��8S+hW	�$�5�	�	$��aK2l��f�
E]Ba�L�E2��D^"lI�m�k.c[��K�-ɰ�{�el+���%�yￌme�0�$�6�a���L$&d��2����Dؒ�|�Dƶ2�[�a�����V&*aK2l�����L�-ɰ�g�dl+���%��̕�m�VĄ��d�2#���L�-ɰ�g�dl+���%��,��me�2�$�6�I���L\&d�法2����Dؒ�|FTƶ2q�[�a�Ϻ��V&.aK2l�]��I2q�[�a����V&.aK2l�j���v� v֞`���^�y���<ҁ�Vh��L\fe�2+���%��l��m��oe�l!F��ˬL\&d��\	2����Dؒۜ�Aƶ2q�[�a�sW��V&.aK2ls�:��L�-ɰ͹Ddl+���%�9'��me��Dؒۜ�Eƶ2�e"lI�m�Q#c[��dBG�d�2'�9��2�$�6����L\&d���G2����Dؒۜ�Iƶ2q�[�a�sQ��V&.aK2lsN-�z��L�-ɰ�����p��]���	����e^&.�2q�[�a�s���V&.aK2l��,Gi�<ҁh�L\v�-ĶBI>��|����˼L\�e�2�$�6�2�фy�����[�me�2/���%�9���me�2�$�6��ф �i�[�mO���Vf�,Ȭ���%�9g��me�2�T�v���S7�&�5��W��(���b2&�/t^����v%�B6ٕ(y�W���Ҹe!W�J����+Q2[�D�f�����@Y������Z=5S�{w/}Mcz����o��nR�B��0^z��Z�xzd�f!�Z�/��s-H��^<��Z��I^��'/>~y�Z��w��Ga-�֋�)������7x��i�`�:�R�K�"\sыcg�s<B��3�M�Q��ju�c���v��sZ�B���\I��KʧC��Z�)N��ԪƵ��ƒ���]�q)B�Km���h��]L��H�U޴�r!X��Q�'=�~�P0
.B��E(�R�b/�ӊPĺ����!F�zbU ���5=0T3���qI����^
A��Kv)B���l�(M:�P�rq��&�5�Qu����E��v{5���1Q4����"����N&YE�wʱn��2�hB��0c.s)B�p�ئ��ہ����} ���-)jFK��xY��P.��d��:�fL�Q7�����FnҾ��2�"��\Ɔ\��Q�_N9��޵NM���~2�7�e.E(���b�B�e����*x�;�0��2�"��ud��6�ѱ����vQ��k�6�-�����JP.�Q�vktP���} ��&uV1z���8tuT�r��&�C��;��/�5=d��|�n��K�E.��]��U�!ͺ���RJ� �g�Mc��Q�eߝ����`����M�㱥J�0}þ7L�[�r�K0��q�Z��]7��͠(9�A�Q�E.\�F�bڦ˭qR}t�U6��]�@wKP.r��9��,�psO�z�$�Z�l��-��"��K���[cԌ2�2t��ƶ]���-5�\��0%��GM˽ZZn�f�0=����)A�<��7=��_��Q�n�W7?�ٺ\�P.�%��w<����co�X��g�Bl'n��K�E.�Y��eY2<�t��M��]C��M&R�̥�rԇ)��,��4q(m�V�X
m���r������(3t��Ww7�N#5����/h�%(�\����<�o>>v�����/��_��ݥO���}~���i�h�C��v3 F ��l�h73aڭ�A��v�F ��$�h��	azZ�H$N�q��m�	7
�i	�	��o���4�L�	&�(��es'��L�QHO�N070G!=m5�p�qp�������vT`8�t��t�����	����(��](N070G!=����0�0G!�̲0N���T
L�-L�QH9(�L�-L�QH9�$�L�-L�QH9�!�L�L�QH9��L�L�QH9��nN7)�q�qRδ��q�qR����q�qR�$[��鸇�8
)g��q�鸇�8
)gJ�q­n�7a:�a:�B�-`�`:�a:�B�`�`:`:�B�'�a�`:`:������,�uwH�J"\I����2;�Q�v��J"\�f���
��W�7�L{hT�]%��W��D�:K���W��� ���A, ��D��EĮ��zHp%�z3ˬ�F�U�+�p՛YV=4*Ю\I����2�Q�v��J"\�`��@&�aK2l��f�
E]Ba�L�E2��D^"lI�m�k.c[��K�-ɰ�{�el+���%�yￌme�0�$�6�a���L$&d��2����Dؒ�|�Dƶ2�[�a�����V&*aK2l�����L�-ɰ�g�dl+���%��̕�m�VĄ��d�2#���L�-ɰ�g�dl+���%��,��me�2�$�6�I���L\&d�法2����Dؒ�|FTƶ2q�[�a�Ϻ��V&.aK2l�]��I2q�[�a����V&.aK2l�j���e"lI�m>.c[�݊B�e�2+�Y��L�-ɰ�g�el+���%�9ǀ�me�2�$�6�J���L\&d��2����Dؒۜ�Bƶ2q�[�a�sp�����e"lI�m�%"c[��L�-ɰ�9Qdl+���%�9���me�2�$�6稑���I2��d2q���˜L\&d��A2����Dؒۜ�Hƶ2q�[�a�s8��V&.aK2ls.*���e"lI�mΩ%b[/���%�97��me�2�$�6�8���L\&d��\m2����DؒۜsNƶ2q�[�a�s���V(ˇP������e^&.aK2ls.C���e"lI�m��(c[��L�-ɰ͹%el+���%�9G��m�L\&d��\�2����Dؒۜ�Tƶ2q�[*c��j�C�Ҏ��+�d���t1��:�DY�M�e!��J��<�+Q2o�DYȕ�e!��J��|�+Q2H�DY�����@΋�ޥ�������ҫU��`<x��ka0>���е0/^z�Z�c�x�-�ka0^��.ȵ0/^z��Z�/��pm���⥷����R�x�ug��\��!F����4%=]��`�\lPE(ۓ]$�ke�8)GS��Nj�K�Nd�.ۥ�]�P.ڥ�]L��H�U޴�r!X��Q�'=�~�P0
.B�h�"��v)B�����\T�>Ĩ[O�
��O���j�q�~B��r�\��"��uT�r���P.�Q��:j���Ҩ:�sk�Q\�����ݘ(.�Q��:jl��IVQ�r����5��>�؆�\�P0\.��#{;��)q�&i{K���R�D)^�EE(�{52A[U3&���QrZ�Q#7i�؂�X�r��ؐ�[=*��)gy�л֩�1��O����̥�"�A�ClTh��s>��^o#%�è��\�P.ב�n�ڨF���&cT�E����8���ǂ:*A�\G�ۭ�AQj����Y��}��7���Q	�E.~�4�Z�0������mk��.E(�tZwa�V��4�6�K)q����7��/hGE(�}w���SP�5�F7��ǖ*��8���P0j.B��%�ԏ�8e�����fP��� ��".g�g�m���8�>:�*c�m�.���"��Q�sNVY�构��I^��';�F'[PGE(Z����ƨede�z��m��L[0j.B��/aJ6����{�&��Z�Bazbig�3�R�ry�oz���2-��.�'�n�~H)�u��\�Kt]�x�х���ƱzG�B1��N��)З"��\��>i˲dxd�|���4?�����L��Y����S0\�=YV�i�P�t�"��8��Q��6C?��Qf�X1'��n�Fj\3�IG_ЦKP������n����6��_�ޑ�����!}�|x�i���m���p���okfd������|}�K�O͂�q+��·�2O����.N�Q�Y��Kq�\���V�ڵ�t����x������;+ު� [�h�[g�y��t�/�w�'�z��<OV�d�Y۪�i1j�J3{?��|_d���w֬�-X�pu��*Ǜ�k��H�����Y�L�S�,W����ɕ
w|�����Q9S���U��j]�X��*+��팳��f��B�5�zѷf�v�Ʌ��5��5�ٟ~r������kƥ&�?�H���wc���ǿa�Ǘn��}|ո��?��xز�ں���_hr�+o�o�C�8�_�[2����?��?�����Mw7�����������Lg��/13�%�z�,��B����5�D���p��Ҏ��[��rʛZ����Ғ/UQB���`��-�|i�rݠA��8|A�dp�¯�=S�t�/l�A�섴~9�_�����<��-7��X8�:�3�]|�g ^�|cI����f��� �����t�\�Ix�1����7ßX�t0�p��5�7V�K��AW����M��ծ��3@/�e�K���@/��3B��e�,��3@��COv�y|�uoD�,��쎨wv�&�zF�{%��%�L�[�r�X�n�8�]���!���`��K0,jw���'�����=1�[c����ޢ�`�$�otbZW\�������c����}�|?M�'l�7�nǫw?�</���IS5�.�A%�j�]�J���c�,�!v��*YTC�R�U����%�dQ�K@\ɢb����E5�.r%�j��ʵ��PO�|�� Z����@C	 ��OY�kyd}�ǸJZ ]��xJ�]� ���z���ܵ<ڹ��:Z���O��ky F���*@m@m�G�b*iķ�)yz-� � Զ�)}{-�����c<%����Z���c<�����W��z���0�� =���N�ͺ��՘S���%@m�1�@m�1�@m�1�@m�1��Զ�y Զ�y Զ�y Զ�y �_j� ��z���z���z���z���z�� =����� <h>�JZ y��` y����d<ܼ�t%-�z@m=@m�1�s �8���-0���z��Jn �����c�W=x ���s���Q��@W�~�������WY��t+�;{8�����Oof/���A��7;uZ�{-�~l?,?���l?������l?�����(l� �����M�/���G`~zӀ�׀��G`~zӂ�ׂ��G`~y�$z ���!�束h£x��C�:3$4ü�mCt4fHh�y�0چ�̐��Ng��Q	�!��m�h�#0CB3�[��6DG'`��f��ãm��P�	�0o�G����a>w���F�)`��f��L�m��S�	�0��@��b_2A�)�t�fHh��`چ�8̐�� ��q
�!��Mh��0CB3̇��6D�)`��f�g�¡���0C=ˉ�����|�!�8̐���C��q
�!������gG�;��0|��,F8�@e��W��R��	��F�8�Xt�fHh��i�06�EG�*-�y�k-�y,:�3$4�|"mCt�fHh��47چ�̐��It��!�!��S�`:t�fHh�9 چ�̐�s���K3`��f�3/�m�^�3$4Ü5mC����t���a�C/̀�a�ց�!:N3$4ÜimCt�fHh�9K
چ�8̐�s���q
�!���4`zt�fHh��7�͒zT�����6ïz5#��_kat��Q�GG1`��f��m��b�	�p��YK�}��,d8¯|������G��g������1�G�8�����ҳ�|g�Ʌ�� �hN����ȣ# 0CB3�i��6DG@`��f�S�]زR9z����:���WZxN����u��^�3$4Ü�mCtfH��|��,�����k��YY~�Zve�yJX]�j�Y*ו�g)XW���_]Y����j�1KU�ֻ��O������[`��R�J��K��~�,M�Z�Z���m-�<����յx���kj�x��� �*;w[S�&�n[�������P��05>�}�֑U�޹��=m�[�Ͽ�o���Ͽ;rm/]���z�����h)��(7�F�C���1��iJz��;�%�-��'�_���N�*��D댧�t�"�^+;�I9�ZոvR��X2v"Ct�v�И��N�n�-��A�?a��4�i�ɴʛ�W.�:�5����O���ʟq���g�QT~n��`�\�iA���N:ׇu��8�J#�����0�ڏCHڝ��U(��{6-4�"��*Ђ���	��ʟ��U)�;Q��M�kJ��L�͸�F�7�jj�wc�h8U���NT���F;�d�)Ǻ�z˘�	a��0�mX���H�?�Y�Α��HӔ��a;��%E�h)�C��i^Q�s�;��������]rZ�Q#��o�;����g�?6��V���r�Y���ujjL7����i�=�������b�Bå�����*x)yFݜ{~Q�s�7�]��X��d�j��U�5cǖ��x��%���?q�4:(JM�^�ݹI�U���}3�Y���?�|?L��[-wCY,��o�����5����ʟy~�u&mUoH��j����s���i��Y�/*��&k{=5X3p�q��x���8�C߰�Y�+)����~L�)k=�w�4�.6����@}��E��<�K��Y�B�t��L���{��Xc��K=�տ��g���sNVY�f9g%i�W�����ɞ�Q�����]��������u6��7f0��1oQ�s��dS�x�i��hB˞�jnΦ'Wv"s��Kʟ�^雞h�L���4pә���!���;�����~t]�'��ȣb�X?���<��N��ќm�E��<?9듶,�p����Is'�54�d"�s�/*N��0��דe��&uMת!��H������?��b�v2���ĕ��S�H�k�>��϶����������y��0�ǫw?_�̑\���*��9Z�!V��r0�C����f��X{�o�m4������6��-���vT����N�m��U�٥��vq{���&�0���%,]}Ϗ.�����%�ɂ%����$�9Pe� p������P����)%��%؃%#�CJC�CJc��%���%���]0�9(P2.9(P2�8(P��U����7��J:��'�^J��C_*��Z �{X�?��.=f)���s�g�+^?�]� 9g�k�Ԭې9�F/�)]M��r��fN�j�9���d�����UEW_bk�lsm�؞��P�L*sjoo�����<��V�5g�,خp���xή�aW�p}�V�$���w0[��3Zҿ�զ��Js2��L�����5�N������-�A
WҪvy��,�A
W��lE�jrI��	a�N�d\`W��V�DX�D6�!K�D�^��d�����,u(����ؼ��q��v*� ��d�	FT˨��u'-�&�{��j��P��J��Z;��W˨jb{���dd��h�&Ԇ5~q(���e��Y��������O����!�<+q�/��W��]�O����~������/��Kf~�>]��K��R�_�O���R�t��_j�.��K���h������2z�e4�i���h�����47?=�����g���(�l�[���Bs�гYhn�l3��y�����|��]̳]��.��.fn�l3��y�����{�~��xn����ۏ�����`7f�o���Z{sh�5v�p���ƨ۶o�V!N9Lc4Gx��K��!'FBSd�M{�g�h��􁱦v
��aG�|�g��<Tr��F��0s�!��o��g�y�����{k\�=�9_����Czx�My���G�����w|��tc�Z���D�ƴ�-�d���� �n�Zn�޻n�Tߺ���Ek�u��~�͐��3�O����ۻ���ݰ*Z�����e�nG�j[Q����>=��o�37��������+��oZogW��^����|��2�����~���y����O����_uE7�Ʋ�_�4��Ʊ5����uKf�U��}�Џ!Q%�F�(5�^+�ۮ�;j�k�L\��wl��uhe���Ҵ�m��w��R�r�ڥ+���k�z�ㇻ��l0������]����|������O����_Y��Ow����_����w�����M����/~L�~���>���קۇĶ|�����cw�i��O�������|���o?����yr���V���a�o�;�-V��%�hln�����Tjې��X\�o����4�p-����-�x���_r����`�M��[�s2�op7�-<]%���#�����R�7Ѵ�K�m_Ҍ�i�?��hn�O�`�~�ġ����Ui�2�k������`�PT?E��򪼎7;[��>j�����o��m%6k,�:���_"������%v��6Fk�i��d�DO���B�ě�>�@�{��i�Q�8��]���'r��&�k������fK&MQ��q\GDj�4)MS�{s�XV=E[���ݚ�:����O�M��'r}��	����������~w7~�e�G��*����"�����w��s-�8&i��V{Ǳ'?9G�v�"mUM�$�G�ױ�6����,�f�o��������=�� �������p{�=Qc�z;$��Q���YC����x�qa���1p��E��*���>�fHe�mKRD��St̾�N�[�v���l����ߞ��O�6���M�	�7\U�4���K�����H���d��e�9��vRC�`�!�Mn��XY�V�u��i�<����1:��e|�׻a��1�~?����/�M�������ؑC{͡<M�ћ^5��x}t��Fюڢ�M�|��ڄ����_��W���wŵ{W\ܿ��?���h��޻b��+�9�|G�� ��Ӷ�����:�|�������+n��ݿB�W�ޕ�}�����n��ݿB�W�ޕݯ~�����Y�k�x���1�ʞ��q�ݴ7��N�>5����F���6�-{;�kw�'�V_�ZG����X���y����ߧ�c>Ly������]/��?f��]��v���~�A��?�O�������<gw�Mϔ�_>�ا�_�~��7����,��{�X�t׬E�?֏�͹i(ϛ�`��֗[�y��4�`��,<N�β$�ȭ��*����f�]�8�d/s�l�|��]f��_����G�m�bgn��=�5�F77��hxx��^Ŀ��ޗ���Q�οO\���_�;}cB�82����ؽ�j�9^�蛖Dܻ�H�{�$;�������9��7���`���i؉�s�9֍���8q��2'��ŉw����_N��_��r�NL7�5��ۓgъ8qс�2'v���CϿ�s����KX���S�ܸ�c���G��趓~l���3� k�-�����.���Lj�t�'	��n���8E'bK&vL<�!i�Ӭ����/���~��,�)��Ӎ���ްhhӆ���WVf���tu�.���2����i㯿�^����7��Ϭ����l�Mޡ�ɰ��	�X���=�&4�c53�kU���kb>�l�����ȃ�N����ɣk�￺�u(�����	�n(j)F��xM�u�r��uHv��5����� ]'O�lw���k��Ѕ܍�=X��d��w�sv����x��7sth��'g��Q��8NQR����^�d����|U������:o���(J@S���ˋs|���co���_��)�9T�#�P@�v2؍b�oj�;g���w2����<S%;��K/�k/#�$�XH�˹����`�5��q���b�N��m^��kow��P$�Ϫ�2�LQ�r�p�
��n�h�H�7�&��SI�l���:����4�0N� ���G�*L,��h���!�£}%����*���`�۶i7S�߸�Sr����E�峯��������=�Ba*�S�;��/����D/_�����G5���_f��z��'��i����?<��ǿ��m��?�Ƿ��?�6���ջ���MZ7黫�︭u����ݸ���T�[�t7��*KI��z�~�#���އ�ۻ�?t�?l�~������O���U����w��w{I?���z�I��z{�����k{���M�����C�FC��7�7���:�h�*}v���=�h�+n;8E��B��N�5�qP�g\�:1'ڧ�y���]�d�-�/U��f�暓�Y���nS�@����:�}����	�=N�y��vS�{����ێ��讹���yjs�b�ɬr&w�s���ҹ��>fA���Zr����J]��[�M,�Z����k���;v�Ytҵ:����D����PW
�U�r���+�uN�]�:G#߃TJ{^\}PmV��\�^���Bv�:�8ȡ�R�q�M�t�8�Z��q�R�C�(�z���
t�StW:�67�KE��t�E�GJos~�?,���Ŧ)ym�.FESD�i��.E�]�u�*]H/D��Y�m�s�`0S�1Z5�Y�UH�^9�9�]�Uv��͹�����J]l�~�9E�	P�{)�3BM���`�vȹ�)�۞������/�ڔ���,�C�\��r��je��SrW�/'��������]�H$^��1[�y��*�b�\�%s���#�)�o��碋��T�y�VO�];7@z�*{z5��U�Vw_T�}Q��ԩ���t��*{YV\���
�Hq9Aw���qU~N�{X���L���椧n�(�I�+{唘����Vp�W����Kr�C�9׋�������Jn*��Ҥ��>V��0\��]j5T��^�y�Ѓ�B4��C�*��09��}�y�O�p��7��������r��zO�N�{�mp�xzP?���^�֏������c/~ܫx�G�Qv�^Й����o���� �T��7q���֑�u�,ȡ�v����#E=��{�捘���p�G^����z�ߗ�,�֐]�2�3��t�3[�<9Z��e����9���h������)%kюwn�zm]^�
�sh�{�V��;�$>��ۘn�tr�p��|�m�n��4�G�rm��ػ��.�����J�;����xj�G�%�yx�id���������/��^�
c��E9�3�v�5nw�9k���2͂��b�m+�e���@wi�܅Z��4�q�K���ϧP���^s[���]έʮ��V�]<�]�׸K�w9�˸�Q��bj�mo�.�.F�]�G�V4�z����������2K{���V�܌�֩�y�z�y�j���N�}|��)�NgN|G��ªjN�p�������m���ջ��n�w����Խ�����=�?f�g���p�?�����qx�����o�PK   ��Xyɜ��  �  /   images/110f4c69-ce42-4daf-8800-65b9db14e3fe.png�y�3���tQ����F���E'Z!����� !8D/�[⢝Nѻ��{��|g޿��wgv��}vv�_vgg6�P_�����DKS�:��� ��bJ*�����K�����������I:_5sߗ�N��0(F@@����[���^PAO�s��=c����q���W�AO�]{����s�|ǋ5���5$��/�}�6�av�B��0��Ѷ���*��� �mik��Tr���ArlIڥ�z�!��lS�I_������i�|�J��?��!�����"L�L�f�>M�8�~SP��v"p�_��b��*�i��:�����X*������#�F&~x������NG�2Jr3��?�P�sH�{�>7��<X�̠��A8po���k	l�ʸ�x�cu�����[o�Y|��r��q~>௳ .��P�m�^��H������e�/�����$��4i�80�o���j��C��ޒ�<�M0Н7!���[v\T���D��As  ����؎>��8;E*F�Z'�"�o��x+�G���Ǫ���8�i*7ls���Ef�;��&�f�o.)j(kX��㉉�4��`=M�¬�x�W��Z�Qj�5��.'%lNVi�����ZᏱZ>�O�.��鶭LP4�0��F�}�P{�����m�9��#e�I�NRۯї&G���k���ֈ�h�54�
��ܳ�=ӄNzۆI�<��ΰ �8�Ż&���B�/h�;ykm�|���ks�_T4�-:���Zt]:�U�QL��X�d�M�P"{L��<�8t=�º#�QR����{B�hh�-��j�>�
�V=��d����~�?}���Ԉ��˽���[PUS��H���,WkD |��k]��!��8ex�y!}:f� �TP�#�x��(�l��e.��9�.�G����qy���{�0�8�����y�VN� �t<x;:[_��E׫���O/(�����C ��/�D%��{�&���R�����Ȏ����l�	��q��9�g��0}�)���$+���<�����?��tl�3j�2�I'����ȭ�7�5zW��=��!HG=o�_��b-R������1ߧ?W�c?�&����l���'u��ٕi����QMrˏ�}�)8!�T�����_����������ƅ �fO����1���dG��
Y�jƁf�?
��"���F���3G����G��e�>2g-%�4����!�c��)��rB�Ƕ� �v��G��%G�a��PD�F�/�	̈́Xbz������?���-(�� O�vA��a�{�nq�iGᅂ�_�"m�j�$^�p!ZVgL���T������Nv[|�}NY��(�mFz�׃u�Ѝצ� >��,���svSBy�:�K����e���vx_�JX���k�|-�[��NZ$>����gR!;g��<��6�
���ei_(l�����9�LV3�֜2Q{�(�~[�蕇�Ld�"�gttE\ݞ���mS��bt;�f�&�P�c@NjB��aa~�y�&�����Q�X�
p���S�L�n\�f�3�E���s���'�쬨t�؛r�O�u�f�֩��	��t��:�Ȼ�V�����-��!:�	�P3Fo���I� ��cd 3�Q>��k54Kl�xg���sI�o	%������lJT�'����:�6Yd�7��e��|t-i"a9u��Z�������#�����_Y��W������P>�ɥ�פ}P�;�_)Tu����O;��Kw

%��,�%��yܔ����nH�ʇ=���Ҫ��p���O��,��Sf�F5��T��NOF��NKv22bh�p!q�ؓ�����I�%R�O��Mw��h;���i����Seͯ;� Hզ���Z��N��W�:iֱ��wy%�7q��>du)��b;a��3�y�0۞*�h�������`��V�}�0~��g�E��&�>�vR�_��=PΆ��W�4hiŦ�W��<�̿*�0��e��Vt����aG���.]Rdİ�p��b�]d����&O��U����@*��r��o��G���}~9͂T�.?�0�y��[�v�xc�>�sc�o;sӉa��1������6"?��[m���%�/��1�Xs:o��%a���2��D�w�~�S.Q[���?�=
�KE����� �$P�"j�8��v<~{dR�����j��l<1�T3�d��%~#�`>ߒ���IҙK�q�l�TS<֯x�po���\���׀l�ʡ��D���
R��A|2�jB<�τRX���� 1Rc��R,�mq���@Y1����ݞ/o�?a��c�2�.Q�t{�D�-k.C[������U��.D�,Z�3��Ge����x�\i�OWZ�	|�#�b�@��^���%�,_t8�|]���t-%�1�y��V�qC����T��žډx?�}Y�[>;*nn?ˌW��̡TO����fOM_l3�eg�K,WddW[�~Q�EZ�����FS��,c���g���ɭ	#�F�c�k���-3�����S!n���T��11v�՚�
�T�����O�480��X���S�]�`�X�RU�6ŘF�&^u�	J��1_)�@��$Ĕc�t�P�^$�%ETZ2�O��E�`�iN?$�֖f\Ծ��n�������Xd�hO����!�=�֊B� �>;�2������&M��4�J�
�4n���d)ЧO[����7]�$��tO28��@<FӦ�,&u�������DӺ��F��*?��#��ٌ�%f}ƚ����G�垛�@��pi(���L����@ӀT����5+�mA�ؗ��"t�RCR�o�1�n�Օ���A��_��ӵ���}i.(��M��`ܖ�	�ʦ�S��N�Ԩ��X@��r�ݨ�+|��mg��&'|�D�����l�LW�h�_ז�+&�`�C��gx�;�H��ӥ�v�~�L���k�x0j��8"��>�����;s��,	�w�ѫ9L�vE;��c���n-M�g�O�#�@�k�r�_�φ��1���w�/�~��N���S�f�u���X��[��N��%�DjK�r��9����� C�R��xtMM�Jfm#^��1/\�n�
�Η�jra�\h�1u�F=��O��9
�ʄ��h���~�>os�߫~�'Fw��D�����}\&eE�Ϳ
B%�ڰgF�F�j4���J7����s��sY3/����]��@)_r�T�Ǧ"�7��+`�R���dǚ�$[Tt�II{�\���Æ��n�n��q�^.�E0G���#��u���"z$1�p�а=��-Tf
�v$�&*VKN��Ɛׯg̋��ʹ�o��b�Y���������:K$��@t���P��E��h�+��,� ��P��z"5R�dEm�^�|����;�Io�G�&T�%7k�rĩs��^���j|!p۫��!�`Dn�f�%D'Ѹ����v�	w�� ��o��r�� FT
���7TTj;�@+	9��c�<ϟl��V�W*��U�����M�F���|o���6�b#���T��htl쮏�����2�`@9���<D�U���+o)�b�r��2pV������D^�O%��.�W]�����V�XDu#la���|k�Mr�����j�sG������P@�g�'#[�D��sWR tO�y���d��
�M�Ϗ��(���$+7�i���DmNß#_ah�o�~��h�c`8%���s��?�X�*���	�6�_~SxX�9>ZD(V�J�
�z�`6d!hN_�0�z_"*�� ��#�僖e��
󜳨���Q���C�k�'k�A�N�m8i�����QAW���V�ҷPH �@�\�Z�����v��a<�,A��T�I	h��߸V�87� �:M��N��͹Ji<|�kމ������sI̺��lE�����h,?�ܗ�Ӓ�m�?��t��a�!w�rJŀ�8��Kt�B�A䇋��x/�j�	L%kb}��/# _�7�օi�*[Z�� ���6����辧���������w�맛ʭ ���K11 G�M��G�2���O�Av���Ozy�8�l�\�z�Z~c4`&Tl���/Hs�^*�5xw��R�т���[Ű�n�-6�e�!�Y����z�a��NͰ�A��&��a��-���ZOR�;0�$n1��-��L��!^�)s��b�4�������Ϥ���`)�9z��k���8��⭍���
M��(��_}�ȅ�/OG;$�]����*>R��s
���1�ثq��(߬�SϿ��|���Q���<�T��dǡN�v���O�xQ���n�Y	cx_��utd������ϑ����|�#nd»�����b����r�Fs����J,�WV�v�������fs������f��n�{z���jꂕ�.񾾘Q"j
Z��d*4Sm"J9�[����>�zӜ2�]�R�S_�|��n�I7M$�{�(�M#��X�����]�T�ک��1�UP/t��&��^P3)�%Σ�~��~Y�.e�I���a���|��h�׉s�,� �̅{T!fg���|<����vC�4^y-����@���#1�1z&L�-ZH�<�x�TŽ�����#^h�����Ogs�;Ӫ�Ѷ}��f �CXmos��7�Jk� ��3u��r_�/gz����@�j��s6/�1��^~s�bٷ߿n1x�ɚH�c���$"����N��r�=�.�mYQ@f�lt,=��z��pm�(�x^�*�q�sG��<�Xϑ^zv'|4�+�[��-5����e[HaZ�E���)�*H1�LXpND~A%}�"�H�.u���]�����([��aT䝌�y,4q�@F�m!���<e �S>�=��c��Ml���p�p��~���Ώ�٧ѽA_���"�:'6h"7��]��>�����)�Y,��!x��E���2D�C |�3�������}3bFꢌ
Y]�p�qJh7gC�ʳL�2J��>2$Qk�7��*����V�݉5��	G\N)����p�rU�/��.,g��t��yM���n������Ȇ�
�kp��T(�MRS����+��jo�z'����"?4]��%��Y��N� �a�����}3İ���p�Nd��]�AH�fԋ��p���T�T�������C��Y��F��e�9Õ-a97�����|���ß�p��#n)y �d"uO��R��g�q��اv�_*�_��J/y�k��+�Y
���H��P��'ݞw%������զ<~qhzqzǋXÒ�j�R/�A�W�۔3�x����Wb#K&W����ښ��#L݌�ԛ1d:0�Ov����l'ں���s���g�eM���{4�?�'��Gڅ|P�%��s���T�_�V+�g�-��4�*�q-�8�{��s~l����R�jv\��y���;럘g��|�XZ���z����Cqfo��+�eG5��ځR���K>�m�Ic����_��P<����~�w}����B77�2&5�{���2SY�ONp��Yp�4����VI8Yd�T��Cq��I��1I�� ���ӭ����m 4�(�J3;Ml��o^� YMz����*~[�1���Y���b<o�wZ%�<Î�o�u�󪴩71��tsmO��$ٲ�U�8����\x�b�cWl<��T"T�����+R��"�]&i<���-a�ŮՕ��U��3���`�`�P��8�\
j6�����o���4���S�.�SƌK0���~��/q�>w
�q��I�@�7�y0=~��X�����i5=�%MI�P^���=��Za=�~�����dk`�Q^��$����ft2#/T��_���ihD�<�����y
[,�������T��o��sm2�b�#_^�l�ݞ���U���=���|���3�&���B�H���ľ���':���j�M�����~����k=�Ĝ�Xkt��������̈́��������a��K��On7�6�ӡZ��:s��D�=���������m�A�R3�{�Ղd@d��"����O�!|JY��6����(}�F՝����C�Q~�2j��z.06��A�o@�$^,������t'��Qw�X�^zY#s�;{t7�y�'��s��H��VʗlHEXJ4�-�O���jO�?P�_!Z�%[T!<z��VQ��.Y79��$��{�٤Ԩ�Ι��K�*�*̖pf^�,= �g^�^�f��̜U"3Ъti���Km�B+�?��8�����3�j*$˧��C�ϰ�y�]�����*�'d�V���h�v�2�h�uY�p���H�B/��Y?-^�i��uf�B�q���*��ƽ��e��Λ�j?�]��nD#�K���d�=�W�L4���1��������td�����3���0m5��XB�$KU*���>^$�֫�2�æ���U���+�߻}k۞���w�~ó�O���Yq٨摆M��|������/b��i����8jL�X�)��0S�;4��6����f��|�D����V��7�Y�؟�kk���&m=��� ���� ��2�T��J��fQ�Blՠg'ٜe?��|gF��%���eo�2�W�$y�^���U��n婎J�d����N���|M��D)4P }���F���u����M�=���� s�LN�#F<�\h.��fY��>/��6����%J�+w����"G:Ӣi����,�Aj5����IO�$P`�o�DZE�:��q%�W����W����bV� ?��m���C�@�f��@����4�Jr�^iSt:�Y�X\+�)�]�s7���&W'�!c�I��^�|>��`oْ�J�S�?NQ-��I|��b�]5.��b�l�D��Y��U�w|�_�D+vE}�u70e&�C�3u�&O��ڙ�1f����5�`Z	�)}������
�u8��io�(P��1{m_	\p��*X�RTX���U��i���z�m7�t�:�5mSy qR�����,n�J��3{�X�Do[��p��6�|�j�P�Z@�8�CpVKL�9@��|i��F�jL+$D�^�݈�0����j�^+�?��1
?Q��<����,]���c���V[��/�!%f����Di��;���o����V/{@O�����e�����:؜	�����Z���?PK   ��{XR�/�+ �/ /   images/12438572-56ec-4fe3-962c-a8f31caef061.pngD{T��vpwwע�ݵE�n��=�w(^��;w)�w�/�{��d�gO��w�yfw�peEDBD  �"'+�
 @�  ��a�Wn1�����_�  ���7��ǿ���RZ�_�̜�Mnnn,���NƆ��,v�����  9@NRL�=�x�͝H}nc�d�𴽱�A�ɓAN6 ��b9����bla�j�~�8� /�M�=-[e�p��l��g��2�FS�Jg�"��c���A���y�cz���(<E0�8��0���>2r�/�yN��:�8���N�!i���<-:�s���\���)��1��w����?� �u���\$><D6f��F5t��;���9�(#�Vn$T�b~�U;�����x�J,���Bt���/(K�i�,�_�ޝE��*I}<��M�|�b��I�۰mʫ�}Vd������1�'�@9RT�}y�0�X@ci�M�(��(t����Nȹ�[$Ǆύ���?����;�2`��.���Q%K{0Ƅ ��Ö/�G�8*�ٜߎ���XT�w�IY�ȗ�"v����O��Nؾ2��a���:�I�G�k�Rx�1�@�	P��X�	�অ!��1X��9! 3��A��p;�$��8�� r�H��z3@���@��b��4'����W|c�\�S��rP���U`X먊|�.?��4��Q�ͳB��}@rO][D�WC�]���G������ݵ�2274����v��_[� �WAs��̔p`��ʭ���j#/��,7
%��A�h�OT�c
������R�6�*�*�u���K	�Q���;	 (U���b@�-���A��f����8�)R��$=��݁���Ħ�뻱�~�DD����:oڻv�&0ҳ��|�[��g�g�Ň �8A�j�!�V�Q�C-[�=ʫ�~��ѻ"����B/��f���u -�x������$Ն���H5ʺT�zl'�i�s�,�ob��X] 	A��g�ontZ"�I�.����vGt��ֲۦ��q����`^* C��(��Vu��(R2Ա��/T�(tb*��8a݈��]#}F�������@<��<y���x�iR؀�ڐZ~������B� Y5|�蒭��|�d_��(��FK˗�D������Ҧ[>�~���*��>5�>X��M���o������+NA�Md�d ��~נWs�i�2n��o/�o���w������9�C�'��������_>�"�f�|
��X��E�A)t�݃�]��г(�3v�6��^�$�G��~p����X�}��?�0���4��$��/��N���J��l�=�b��X�i!�4��`�L��210K��7��o��]�fmD��a<�}�/H�n���eK��awZl��3#��	��ذe��B�9��!��6��5p�p������DQ@�K����
�0a�⌮��N����t�K��Of�0�ߛ9��qv���C��܄OƔ=D0�d>E�)�˅�JƇ#��	��\U7'�H����^��Xsa���w��q��a��i>�6m�Y\u>�S��g)�,����ǯj ��$0h��E�([7�/g��;���V�"SV&(	�9X�EL?�4���ngk�RȽ���u
W�?��md��'m��J��T&���/��B�qg��S�{[��@Z�]y���>�8�Is��v$�j^���=%���-��~i��@�5��)˳c��(0Ko<��.�����~4����+˴�x茢��;��(nJ{�ͽ��Ňe�e%���n��=#xEë��I���]�d�\g�HKC���D���V�:�HX>��p1O��{TK ������(���Cd�F���s���A�+ �)���_��%��ܿ��W�
d�J~�ryz{{R�@o?�s�1�?���}XAc�z�����*	������Q&߻�����3���Xe�Z�'�A�omS�wԯ��ֈ��rF�)|������&y.��lLb�;�4=ue�!e��;z/��dJ�䧁�	,���=����7x7��l�ՓH�3_	p���<F?K �V�CM�������Iu�I��k��qzFg�}Mw���DD�94s�c�;�؏�a����c/4l�5�%�� ܨ���ǩ�z����G_�F�߶Hhuv����ѿM�{����U�dD���gᑕ����C.ޞ�ʲ�Raߥ� �l31b��a�ġ �u��D0�����N�|?cp�T�ź6�$A.���>�tr�r�=о�Wɷ)�0��Ƈl0�D�q������߁6u��y�T���p�w�>�ؙ��m�O����"I]�\#1���U�xI�x5� Y�p��~bw�$(���9�� 7x)�2�����v����������<m�MjG��Эz$-�G�,;d����x���B�p�{�:�)��'��}0���k�?8�8=#csK��+��6���0�㡇7�,�Tѿ�aR�Sa�\���-0���]|e�O���:'�G�-g����o����`�<Q; ."ze��Y��4	ywg%���H�x��gd�)��� d55يio���RW�%|���	$�u����G/vG���S�{|�;�K<����_�cX2��H�� $��+���n�b�'l&_��s�*�����g%��7�z�޿�0��n�K������왔n/|0ܾc]�f+[Q!"��wh�a$?,�_ɺ`5 %&j�<���|W�"�8eMol�Pn�f�4�z���2����knh�!�D��_�/{�>��~�J�� ��D�8������#��$mV�7����C?�a�����O�_�-��d�ɜ��!�fW�.`[�z�_�Ϲ��ޘ�3!��|��l��k�9��>}��z�O?��w�z���4~�Y<��3�������_滒��������p~+p��A&t�h��((��a�3��#�$O�a��H���|��J��Yt�U�sw��1>��j!ɼ��E^4=�%ҏ�Ѿ\�FQ�^7��XZdTi�&p�xOW~q��b�%��n�y���2+	,����a�+���F%;��q>��JicL� �vc��Śln��W2��\��S)f�]�˙���ՙ��2lLdl��~�l�?�(r�.r�g�Y����=���%3�Z僯�I��?Q����G~\�����	��Be<�.��h)��h���蓼���iˌw��;��F+DJ����/��ߩK� !XS���w���m�����/��؂�P��=s���V0�ȴɡ2��4؊�0I�3l���q�DI{G5��U�WY�'-VӐe�bwո=����z�T2��yu&&�ا��sNG����=��Ga��w�k���͑ 4��q�q/������7	v�S��"Z��D��0��XX>�Lg4�R��5�א��ӗj��-^:$�B�g3l����LD���irn� �o{�\�oS��5���v�!ck�6�>4�>�-i��7�<����0�(��/�3x��y����Q�d#."DKPPm$ýSNRKX�7ӏ˵����M�2�6���V��jаҷހ�	��imz�vZ��	�pɿSMԘ�Q1�SS���z�d>>�\.Y�"��T�s0���r�A��~q��{`u���K��:q{�����ߋ!l��&�a��&�8��&����L勵/1xIA�Ƌt/Z��:�	����08��c痌���F�g���vF~-�+�����m4ٌ!�6�G�;nmP�%��X���̶w8����}~A�jN��bw�(q�����i� ���#��Q�z����שּׂ����Ξ�'gg�iEN͜4�JS?���}Uy�I�C�C�7��yc�jb�B��x9���!7(L������Vg��g�Ńp܏ɾT�O;7&��%i1��|m^6�/�y�w���&w,3I�^�Ei��aJ��;�A�dW�K�>�!�[i;�ľx�XpN�ڃ����W8zCs���[��/�P
߻�EJ���6������ Z#-ϫG���>V���Q����
-�ʁ�������=��K�����_�bQ(!O�i�o�h��ivԇ=�(%���|��m-\����<� ��]z9����	�`�i�����o�=��=���ۼ��@ht�`t���8�t��˘���ԔQ�P�cA���VтS\K{�����HQ�������{����=O�����Ū���e�h����݀k�>a"fԙHaUG#��w^y��/jq�/22�DS��&�eP�sfR��0XF�jp��A.]f�=&�0Q��� �"I�Ϩ����a����6I���2��1pșg�#�>q��׷+z�Xl��E+�īӣ|f���\���[2����zX0����?��p5*J��c��%�#��A��]�pJ���B�BXJ��
�E�؟�B!A���?8�����Mg�ݳm�6�^*��'!��mL\�++�/OQ��G\��
т2;O��<w���tB,v&L'�O�"���4ONx�na�v[lq?�}�n{�֕����5��*����3�~�-$�{�5�I.�������W� Ҁ��r��ϿY�8�P��=��g!�j2�(�H�y�-,l��(CC�1�(��aA��� ��=i����q@˞�ai{���x���e[��¥Ow����7`S��:}��|6�fd���Ut��&���?�����eKK�1Bn�a��mWt��L3�'f����CjNYp6��u�Y��3��8����a��/���#0Dz��;�=w�HBJbsz(>����]��l�X��vB����HK��L-���)*�A{-t�x�3�������?��v�%��m�Y�u�^$���8	Ptn�?&�֥�:-ir��ԃ��j;F��U�^J�8!Bو�����u��Wo��\��� h����Zv�}ȁ�7�8N�����T�vT�.֐���K!�b�=x��:6����5ӗ��+��9�>���og��:���`�F��h��� ��X��
�l��b���,����_���䥃$�E�ۻ�n+܉����~|�����i'N�+QW�~|��ܴV[hp^4H{����q��6�ǔ�=$!~��Kw2��!��m{ԝ	�菡��}�e�b�����EM�������Obb{}B|,L��g��a�H���.4�e�}��`]憙E���u����7�
�;����IԪ���07�a9�ui�!�^�=��5�_۱m�����E�4}<�]���M�c/��u��3F�^&��~�"�w4��ƕ�u- ���%#��H_�
&bqH����	YK$=6�7-,6B�����1�5���k۸�^=������	s֍��I
�o��*�Rb�9�k�W%J�~�-�X����D�=m�1����2E�JV�,�����w��14���i0�W��W��=,:���5�h�}7N}�%�{=$ ]�ƏqS�������-l�GB�δ d+i�<�`��G�~�^*����uk��q֝��R.���9���X
v'�U�Qn9���+7�c��C�89�M�UDz��D�6R,X����v�b�H���K_���s;�^/Z�Srs����2�Km���0�k�q�TyX*U�	�5C�\d�|��3c�\b�4�C�]���$�gb�x�-q=R����'��uf:O����P�nP�H(]N<h�u�.�[sgyۜ��M���0Q�>J�Y��ǰ`dq�i�e����P��%#���-�ȏ�����Q\,�
��O�➴b<˹@�3��4"�}LgB�;xB�3
�2:?���
i�[��4�$21��M���W��G��-�f${��W�B[��1�7o7Ľ�'�uCd|��*ݎ;���Ҵ�\�C�gŻ؀^_Iy�"��@���{�;Z_9c���w_��� ��H�GG�V�Yh?=y��,��U5&9k�mőV����ގ��sa�`ӗ�z��~`��@�!c����d����Klq�E,�E�R3GX��X�+�N������Ӌ�mV�j����~;.,�/���N�8�_�'r��m�)`�&���X�G-a�E,��A��Ƒ�G2 o�Y��/�`ڝ�œ���)�؍y�"ox��n�9>��F�s�1a������0�|���S]<>��?��Z�'�l��1a�;���`��(ei�F�C>�ȚVMP`Կ����re?B+&;�m�vg�~<�-��W]$fzm ������x�"L�r���m,	�Hf�
��63�
� D���F/�� 2K50I�������Vn���Ph2j�V�F����������˜&Ҡ�$U���:}��X�ܑ��V��m̾����7G�D,$�+{Ӽ��:]ҳ������Wn%��ߪ۟r5��:c�|��n�顬S���٨�����0uv�����ƻ �㧕[k�O��T�u��W�l��w��͍oi����=2R	?��36ÿg���O�ߚ�B�t���z8���wΒJ].�^�:^���Y��B~f��/�,�SFX�������}�&"�&|�
��f��:Oi���Z��դ�yq�X�r%O������dЭ3����?&���UOj�~AE�͗��h�)?�:D�-�����#r衎c�'1�N��a"s^�g����2)�%
��Ʈ�9�(Z�L̹k�@R2l�[^?=�0��(�&i{ ����y)��wZ�4�#��k.DM�H�jP5���B쯎�͕�*���kD� �n5��u���"�b����a����=-?/�p���<2h���g��!���s��*�ENT�*wd����(	I c;A��/�B���;M�^R�t��ɺ���t������$V1Rϳ��FZ��Z�-���b)S�-tS�׶V����C'�w̝\H��Y�z����N�~�,gլ^��a�1�|HΎ��U��U�~9��h��!f����`d�n�=�C�J�^�5�G��DrF���2��j�hf�D�V.��1P��9�=v�Z�������K�?>��QK1��K���l�s5[غ�������IS[��-��
"{ӆ�y���	7WL��,T�c+���w#F�m8���0f�F�Ҭ���ǁ1��1��0i��R�oe���aFj������:.2���,�p�����^�gTO�Ql�͠�0pA�ڧޫn�N�|?(ڎ*G_t6�����8�R�"���;$�ٗI0���JȜ"��_<.�.��R�r�U�P,����	�?6����ǂ���r&4�Ե���R�N噇�֩.T/	�U���kl�~|�Q]�N�L����ו��G��y����{d�!���X.zd�
�P+�e�[�����g�!��L��_|MuX7L���Ǒ��O���2�^n�����w��Q�~�6��PF���������-�O�
r�t�xu\9rB}��^���U��ȱa�Y_
���>��si�=�"���D�c�h�Xt��T�ƅ���[�8	������Ҋ�
nۋ1�d�U�jS�Wsiڣ8�R���h�՗�|]JI�σ�����K�>�ƽ�壠�6z�T�ocG���o���>(T�o����
L�$T�1b���>�	���e�Rn�呾D�hh�2��E�)�r�Ö���
�����Ӯ�}�����������S+��
�=��e¸��n���J��H����&��ԅ�ڗ[�粡E}^]N���rP}�ܝwm;4���%�ٸ���k
�J${i@*�଱�o����Vd��aB���<t����!��Ƹ�j�R�]�\b��c��&xԯ�{_�º�w!pw[=`��;�\�Lj�}��7�d� D��`��Y�h������U5N�W�z���ב%�������e�ud�10� #b���	���6��	֏�j�����j�O��b�U���iF��@������@^8�P�}%�h�֫���5�h�6A'm/%y=�o6��B*&q���^�o^M��y��[�� �3�(��C�H�B�ܚ�[��/���)���XjHST������?�s"�xI�6��l��)��;�y���̬��!ve����(��O�C��ƻwăS��ΰ�&�~�3� u��o5<�������U��\������2$���?^f�.�@�j��nPP���&�^�;e|c���FT�C�Lc��?��,�q���}�~��-o���:րY���}w#G����F.�I�ܢ��X_�>�������;私�|�ⁱ�W����]޶n��Sh��؞�USR���R	�JF���kVvoB��ϑ������q~�m�/��bsoMM�n��m���0���9�O+h=�Dc(s���3"�y����R0#��j�?o�ʗ��q c.*����>��k>�B���;Jsj��K���hEޕ�>	�l���� t�n�7���"���ܢS
�z��>&��n�k��-�U��3�*���c}Kĭ�Y�#�����j�͗%z.Jv: ���8o�6������jڏ����T���>��d�l.Vwڅ�;Dc�w�__5��fe�X�0�ht����������1@�c�,�����8��F�]h�9�����[i_�.<ߘb3�g�TU���8��W�`�;,��
��r��Qp"�)������Q�ئ�fS�	�84�( ����Rd�М��`7��#;�U���kHS�O; c ^jah3��6����B �k�Y\R疗K����7����8�cH�e|>��׶�Ț[�z��Ǭ���R���m�.%�n�}m�vEs%�V�H�s[]-"��%�u���չMEs%�OD�e����eŨ�΄�Wc>�J��кdFfi�m%{Uh��$b��jjXh�������b.�,q���x�e��)4�'n�����^���I���8�zpI@)�Ͼd���ݔ�Դʘ����v��"�g������K����M=�
���2�j�7����Δ(3�_#����F�,�z,��n�qh{��y�GAm�;5�n�C ��!�Ēϟu�޼MY��x�����7�ٵ�eb�J�vr�Z
����@�\̋�6�Y8�i��4����N龀b���YIbo��>=���Ȳ��Qu����DrS��\������<�`��봡��d�o����<n	���.��̇��^��H�����#��/�W8b�W���m�jb����q�����I�Ax%��&��6Xsp+Kd6`�Q���y�GvF&����Q���3.�a��@2Q�T����bo4r/
�7����������z��@�"��2 M�9}�l!�鲥�������Ε���ʷm9�/]@�XϢ��-*#"ZI/�����
a��5Y����GB�3��ҚK��A~�}@\<���^�B�[K{�����R�����)!K�N[V-�0]02:fͬ���)���GQ�jG�e�T�/ӛ@�璫���/sK]�}�vn.H�����H5�].t;XX�mN&�Ѯ�cι2�Q>��N�'����y0$,�nR�C��M��]N�6	N�`�Her-�=d����vx���c���t�Ʀ@D^��=�a�cU���� ~nA��#�b)��']�Q���Q��K�8.���d����e�Ua����u�yt��k*DK�:�(S�(u��d_�n�y�Mx���L�n(3�a��W^/yr��� ��uG��<T%p-�/|'7�*3-�왓n��Vn���Ƌ�
�$)-�,L���F�^���n�K�?g��q��D��ϼ�<R������@��}3G�[��g�+��x[�"�Z�n�E�Q���EzD��EI��J�$��2xIGId]<]�`�e֕I�tq�hQ�W��( ��4`�tHF?�T"��p�?�@��Y
���3$H��7���U�_K��t02RB>-��iD��E�ڐ��r��Ҳ�C��������A��:M�$k��u�Ib8VWH��$�_*"����[���k�`�V�!K��H͐Ѯ�n���)T���w|�`�I�	$�i�(�H�vYC'ǥ6��\��Y꥙h#�R=$���� ��֚�0����,��Wl���Z��y?z���o+qp�� ͝v����7i��<�0lj���x�M[w���O�l��ץg�̂@�+��L��^�6.g�]xD:``�:�F��8�Z�'v�g�(H}^_�������@�����C	�ܞ�ћ����Ve'�}xeOZ��k-��(^�<~�<D�*_��c"I�%��pa�}�By�����q���N��Νc<����?ѐ)��D��������A���P��m���w��K��esy-���R>|p�V�@��n�)~@BT�L/;�R.�ښ�6X$f:}�  ��u�)`΂MH�-X�A%���Ue�W�G��8�_\��P�'��r���"V���X3"���Li�N�a�K.֗���H��47/�-7�C�w/_�<-j�8��U����1I[Oz s��(@=�]�Bh�%q����{�Y���a\_�  �OFt��c�2{"6(x�4��3����2�^��S�L]�!��v�B��I(�H��[~��(А�Q
�D��5�b����oM1�|��mmIgl��uK�ϩ4U�D�C�9NUd�t,CQM�ok\Hm�T�Q�A2#p��0��f(�Զ�vk�ٺN���O���p�q|����
t�/��2�p��n�tug[��W�n��o��2-�3��.r��2m���������l~Cpnh�Gl�*\�ˋ*s�,���#|r�<4�e�L��Ѫy�Lz\I����׋����_y0~~v�����I������z���a�C�U���d(�?��G�gA��ø��|��:5]U��s7�B��,��iz�bI&ͳ��v��/�&�É�,0oi\ެ^^~��f7'��[�:�lC�f��)��e��������-�.2Zʩe��v�p��<�K��D*�B�[z��BJv�:���P��j,���~�}�ߋ���gv����&!}�u�j-?<)����0�(1)Rԩ�9V����J���	�X���)V�,%�X��dm����a���`2����?�]����ˀ��]�'��ߐ{EY��(4�����V�/���#G�uk�e�z(y�v:p����y���(=��؁L��>�6>� g��Q7Op���U�������,
��ZG�\r�ȹɊ�3u5��'
p�'�h����S��Md O�M���#��:y�I�t5-~| �����,Y����s,}�M�4E��P<J^A�F��`G�SFU�̅ɬ�(I����N��v7��m�8U:���Ę\����2L_;J�����N�F��ķԹ 5�'��U�(>c*�ЋsR�%���~f��s�w�`l����:�P�_`���꟔�l��X���h�q���p�������*)��z�@�N�FQV����@�lcJFJΈ$i����@>~#��w&`�y���J$��D�;�(��!���W���D�J���4:-,�R���گȱ�~����c�On�����dC��"�^8R(Y����9Z�ҢG���+����A�˃z�q�\	W*zJW]eWߦC��+�iddB�S�:��ؾ{n^��Ѩ�WA(pyloNJ}۹�p��pǣ���3ȿ��%RM(�.�v [��N1����p��f ��7ğ��C4�����[K��0�T��uH���=���L��S®�t���p�g���/f�s�دH(!�bTC��V}�j�P��d�;���L���z��On�VY5O#&2�J���`��T��Fvi$n������|_�-�Ǐ[5�!�l�&����h���#�/寭U��l�DL��LXy�"�d��V�Q���S�=A`�cڴ��'՞ȅP��-�VL�N�����M��>m<I ���jFzn��'��[���RS|�b��2���ۚ䌲�f	8�mw~mф=����pi��R@��3�5Ԍ1���_L:�&^?�.�0�H`J�cL>I���G�֠��w[@_��'Zq.�W�/�c�bMg��繼 ���.����ra8��͹�C)Go��%�@l9��YgA�UI�]�?��\�It���͹�n����%ؘ0�+5,�Y�ڼ�g�	���q��[%��6���d��b�I���$�|z�D���]�4�A�A3�ٗ���ϺE�}�>��z��ؤ$`(?a�����p:L�>����)��i �4R��-����(�Jb���Z(4	���/��+��K�����=��Ŀ#���Q���C�޵BD�k�8_K7�Sp�bY*����]ؾ�E�F"����A.�_P(O���n�j�&�_�=� GҢz�co����F,����������̋;���m�Ђ��@��r���ky���n�{�>Y34&B�����SJNN��M�I�V�΋��*r{a�R_�?�����b����6T��ȱP���Dw���I~hJ{��XI'*LfXjmd�FB���\��rf��2ub=v/=z��O� � �R�fG�BB�h�v̟^c��N��< ��t��i.���Rٝ��O���'@��3��/��Y� O&�����ٔWz��[�l�
��|������w����	D9i�}�>:R����)�>(1�<�b��kR8�&Tc��@���t-�"l��-,���2��b��;���i c�m�".�5���h����$)Nl�Ʃ�<C�n*�	;���W�^�՚���֋�8�����N�#t�����u�
U5�7~:����k��#հ�������l�ޡ��u�)+ރJƌ>�t��^�>����L�22cj,1�"BR9y`e���SU��.�b�kWX���X4�Qc�2`IP`I���}�&��`&�#��&����T�k��bv6��}���ՑL�����1��AB���Y��ݜX�d>�Į��ǿ���H��#f�B�n`x%�xdZ�qOg�#
L�@����,p0��7}Tq��0�oϗ�<Fs�P��Z�2�a	����J�=g�y���bzo�,&�a�g�a�H��9�ӯm*�	� q��u��Z�Ǥ Hjѽ^tY-
��U)]d#&)��C�iA� FQȘm ���QC�EC���$�c���T�}���F'�L�%���	� kg������q��k���b�GQ"����?[�|���$,����<M����Y���du�nz�$�=wB�c@�1X�a_�	���7�ם�N����%;vMl�5^7��t����#ډ1���f}��XG�e;�\2HD�و<�«�z'tS6Ӽ��¶%3�O���n��+&��ds�:�g��H��f�P]���4��*������Krz�oϓx��ƞ�)�BO�3�����g����h�]�6? Љy��R<�(�'',����Z�{�^�ƿr7K�*�G&�@и�5���%6:��;E��� ���x�E�h.�m3>e<�=�P�x�II�N=݅"F��[`��LXe������vI<�8E(��l5tl��S%b����4,�=���>16��y�E��awc�'�jf���G#0����o�f�_�GU�F?�7_�x�dEi�V�mG0���'ki/&���*o�^�Vr�j�M�"UoA�鏫����p�yb�%JM
냄�rB�����$���ї�XdU����c#����ٹ�D1�{�S�KǒF��+�<��k��#�ƽ��W���!���Z&�j�A�e5�)���1Pُ�m/5�4������Јz�nPT�������Q���h�m�D����8����P��o�.~*׀;mz�+�w�[�2af�p�й�>��$h��X ���;^>epSo�a^
 `�m�����	�3�_jl9�M^n��C˺��E������e>�Gi�ʧ#�r���r��f���v|�>�#�d�p�Ɠ_岒������
��;��7�g4����HU����lC������7j�՝Lqo~#�x�Ryُ�����K�B�i�h����͋�Q<�u�+\4�`�;>�[�v�b%⋠��
�o��+l����z(M�k���X� .7e�k;i��!�� �,�}w���*�M�I/|Ƹ�U?���p-�X���ئ'D059";~8�	~�2�1��z	T�����AG����M`�ڈ�;��8˖ʯ�&Ͽnx~�����2f�.>�|8�n3�6���s(����{$q��u���o��;=1��w?��*�0�0h2�)�E^ �b���e�6-i�@U��m-��Gƨ�hW�{T\=W������5n;�=�`�n���W���`�{.�3?~�Od�� ��ȉ��Gšo�j�!=�g!_�Z�����vyЫP��|���A�PQ]7:�/�n)���Οu:�Ë%_�]QN��$E��`.�|P���e�������/F�+B�Ji�D��V�����Ĉ�y��i�_��l���]���O��Gz�V�����f�1R�H��a���Ȯ]s��ͻv��hqq<-.�w�#�o51��H�-�x�(�7'�U��H`m���s�s�dؑy���e	�?���f��cJ�Dz�]����c����S6�S��vș�8���S��<��J#�jl��}W}	[oS��j܎(Ñ����G�+�Ƀ��x�1c#��|j
�]�B�\�/��\��B��3yV��.��P�"���d�hbϢ雴Q��녈�O��Kv���äu  ��\�>a`��]�פ�2���~  ^\Ը����@q�f%�MwEfT�2I=	�X�XٜwP ظǒ}��2�	�#��jd��A�U�����\ǊvT'3o�44������| �B4�{���ut"oD*��c3|�%%���~@�F�c���Q��/�~z!�RX%���E-�<�g�p��v��.�������?n�O재ܵ�^ZC���Ќ�W��;gdf��_2a�	�p�\���I����Co�{�ڎ@�+�iU���=j����'��3���2������� um�C�ѣN��Fu���%��҂�K<������bԓ`d�Z�`
F�5��LX��q���qA��sW2���޵LOΌ!�w7!BO�ǎ^��I���]�$�^IR�S����������ؙ��M!�s�'É0#���g��ݒ��ɹ�����j��V4t)�G�� 6����A�9}nC��Li�3�A��7�Ńxj5��\f����,=I	F�U!��I�d��g74r�_�%��*�����B&W�$|j혒���70:�\�;���a��n6%o�|�^��`�e�5}U���W��ל�ߘPr�{�-�V�l�O Υ|`2�ا���f��)�n)C[��S ��1Z��K����(�v��h3�1������\��e�e�BS�J�/�����A�qYo��)��J��&�����s�־'ᆹ<�4��)��R79�"������	�Z_�d�%��g��bS��W��>���gm6�fqHA*�H(��
�űd(���@b��n/��U���$���l0�=�a"W�ν?x	�B�>���9j�D��Ick�[EI�$�9��ec���DL��9ߎ�?�]n�|2�-z��
��;-C��|����ߌג{����p��Gq�
�L����%!�=uQ"�k9p��˲r�i�N�r_tjd����٥Т򃘓�M����.��F5D�out�]t��8��<Ԙ�����z���{p��ah�@�LB����Kяk:����U��~ÁN9��J0l&���T{� <\Q�#�(���/1��#��+!�=�D��f�m���T��w��,0Zn�H/�R!�RqvQ�\������8�� ����Jy푽jb�� �O(�6&]!���7�X_�*���EN#rq �/B_��8����]�<�%d��j���$�����p��VM<
iX.���l_�����n+E�5Ș�}RH�۞�|i�����H��@f�ȇ�sm3P>+�"( �mU:bL��0p�gJ_�	Vq�}��#��t&�Lh��gy��	�]�ܼ?�K��u��by�&g���#����+�I!�]�LV�'>���Ti�E����=��o����#��d¤#<�)��>C#K�f��M����}���XKd�'Ao�I�۸��+Q���#�NQh�&k� �h���|e�#M�`Q�r]�����:�s��YKGT $�[=��|)}E8\�����@}0��E*�S	J�p#��>���w������� �=�O��ژ��ӗ�H��c�sI��f(W�6LAf�r��� �^���$�����dr�-�v�J��3�^L�(8tbՌ�k�S�Qc�&�cԍM~U�6�3[Ҋ�'�Kk��X.'��x��=v2ւk��,�H� Z���k��wf��谮q;:d�7�~�Y��Jֳ�ؚR���oN�Ϗn+���/��� ��l6Z�}�L\�6�_��
~�؈[ڔ-��3s���W��E*������l�r�+E��>L~���;e����+�↶vq���Nq/����Nqw��R\(��Z��Ŋ����>O��0$�K^�YQJ����
�Aq�4�We�p�%�0{�ω��	T]����vۅUh���z��(���f�k��pK%�ۏ�.�J f��Ĕߎ�ͿAP}�X���Y�w�#�^ы�E��J2[v֝6���mʝNKZ�*4T���_!D=1*}"�a��Ƹ�����N-t
Fv:�R<�?��ֱ��.4��,d����6���߽
G,X-�w6ݸ���+7UY���W�^6YSMy�u�n�Lq���I��EYGa�D@]��l�gfb$� Xu8�)d���l�vUkDGQJ�w��6��Eg�VRW�0����ϋy-]<G���GQ��姨�oZ����[���#���� ���M5��� �}x6����5� ù,���x�b���t���.C�R	G�P��S�q�%�_�^������p�un}�:�_�����6�@�� .�lڧ ����,�*���+Aݟ��ߠz+l��o���gk�#�L��}iO��c\\�Ԗ�F3(���0xY0�$Q0/u[�y&.��a <����C~&�zI-�����+���N���7��hÐRzMZ宋☛�;$�܉�?y����T�g����۾�N�k�Rvݮ݁�Bj�;ue�n�0�:��W�:�Ŗ}�״����l��"L����x�v��=\c�w���!����d�G��]�ڍ+�!%�gs���y����m��:k�1=g��Şj�$n?)!��3��:��A�7݆r��#J2T�9��A]J�2���X[t� �5�bQ���ua<�)�Kj���y��n���6��M��S]�#���r^�j�$yB>?���O�?���8������I�~Ҳ�IHf���e��0/�哢Ѯ{ff�P�ިMD���j5�!�"~��Fi�?���JOc�چn�Bɪ�B���i��kji��8Q��Ah�)�'���(@��������2c�׎�ݭ��G����ä$��>/�D�i��GEص�1w�����|��j���f������V���><QLB�1����\�Ѯ�c�G�dDJ����A���!r�:uPm{0��\����2����5��a��؃%'T��˹2B�B*mx�ޥc��.-��7���H����
s�˲#�Z�.��S".x#}	�i����Xp9�[�u��Pַ�Y��@t�4�P�!l*U3i�ɼ6��`_W��`ͻ��l���k٣�	󠥉[������>��w}���l5�e�pP`���"�q��B_w�uJ6)>t]������j�����nk���:c�``I�53���y2(X�mR�!kI;��ċ��l��q�)i�Qo�w�r����{��-	}�ʋY����v����Yvx^�����Ǖ�a�󕓟�ewGjk^W%��[
	 P��EH5��d�-�;W�G�9pд���#�<Z��m��R
/�g+���,��;C�	9��0�����5G <���4��S\�!���S.���Z�̂̓�ʠ��o=��ҡ���R�|؅aH�2�|�$��_k#�V{3�'s]�qǒ�x���c�1�?K���t�>�5��_�V)aϜ�=L�jq�����>��u/HBy��=���P�>�Dd;d5Gn�;z�.���isƜ9�J�=1f'��U�rB񄝆S*6��TdЫ~A췏ơ+{H�\������$ ym�X�Ȋ�7Sn���Z?]	v��V��hw�zE�\7U�a����Y7�������+�@��P�>"'4��؋%��� !p���>�H��,6s�`�q�C,0>�"��!/���l�4b xs�h�c=�썴^s���X�=%	���Ȣ?h���K����.��R�Y��n
�d�sK<DC��5���ھ���^��έ�D���_�Q�ίx+�=ՐN����Y�G�Y>���uZ�W��Y�}�mݾ��?�w��p��,�Z�^����ܶ[S_�[<�w�N�ff�����B1d����:���C���2��{��䦇o��'����Z�r�Zǜ�&&�ɮO�V�l������p����RJ��oU(�JŎ��yfY�X�gm;�"~�7��N*����,�T!��X��;��F�+v/������9��#?q[?/��{lD����o��?�౴���W�ִ[�|���d�)�~�{w����w!sFw�̆3�4����ԲR�`���*
;�,���X��ܵ"��m&d�:t�2c(T�	:� _�Ag�_K���W�D�'�'�.�D����E�l�G�^��x��~�vq��Rc��ohF_U����0<B��Xb.���0��
��X)2�˪�a" ]K>q�,��9�	F9�og!	z��	
P���]s�i�A��|N�1%��46�RL����#g9��%:��[!z'��coNS,+9Q �L����òi���(l#{1~-.(�P��y>>B�}"�#P���6���Ӌ�7<�덷Dll��NAA��P]�I�,�NY��}�.wc2\��E�!�>|k��v	g��_���"����kuK��X��C�G�<���M�q��l�Tz0�1`���L��<��B���/z�~�h�~2:~-��X ��:�a;v����j���wL(���%�23��ϲ��yZ��cT�Q��:/||/Racݧ��їb3�.?�A7�I��)��@[r�,
n�	�=�"?VpR/<�n@䉩��D�����7=f|��1�Q�_rmA��x�T}��F����ӂ/J BJjc�����\�;��n�
ȹ���������d�R��U���,����67-�)m�DW�7K�tM�Q��;u(a�eb7׎�y�I;O[6f�U���	�;d&B(Q)c�i|<d�����6�����IWgqY2����І��˕���:#'I�h\��I��:��xI��3\��-��_����imo�(b�hE�`Oy�㡃jц�����K���N��v�R��2E��ޓ��|Lp_�n�c]��7�bp��Q���5��G=���]�>���q�,����+{�W�O��Y(+W�Ge�Y���c���+Ne�'
~�Z���ru~��wK�[t��!�3CR:6$122.�(�!��"h�.R[ƏU��[+���{��),n=߹�]�Ʌ�L����ʩ�6dɯr�b��m_�TΖ6*C#+8�k�ި�Će�� ݸc�PzU�����X�p�"�&{�T����bkԹ��� T49�}��ا���?��}�+�K$\�"�Itg,�#�L�/N��v���0�fc)�h)������I���������}{ޗN��,3sb�ݪ�񰝞��+d/�vZ(ެ�+dC�����cU�ܙ3��j6�n��)�VV:��R�]� ��~(dZ���f�.����۪O�����w�c�7��!HPd�&�v:��P��m�f��R�^��]�Cf|6ܿ�F�#ސ"����lTFa����%���9[�~Ҵ,Xon6���,:D��e�K{�#�j�09�R뜓�D���t+�{���?�дZ�U�����<���CW𾷒�\��ٷ��]Tn63t�7��܋�LʓF��!5"�DB�-5�֐�a�0�f$M�_�*)��Vs�=�<9C���m+�1�[�������w�h�=C�C�f�
4����N��#�	��b"w~ht��x��Hi�6V�r�|�4�O$3M6���c�p|� ��@ �z�f�z6u0D�V�FĜ��渳����|m�X/�ӐKG��"���4�8��W��Gi���FO�]0o%��}N����ֶ	�Dt���Y�EW�ڙ����:�������Şw��}��~�A�K�������qK�)g���j�L%|��.���Q��v�;�T�G2B�Yh����:ߠ/�����p)�%��U�U�ɢ��$.�L4�w �~[ǆ���>x��״H�`n�3�{x��>9`6{�ӟj#;�+;�d�"����FH��9�ۺE�Q[#�m�WŬѷUr��ǍUZ�Ә�	�5� =/�~���tY�q����~� ��+D�*59������|C	[���PN�P�{o���⮘��g+I�_H������m��=b�%&��p<V�	$��;q�g�جH�O��6�el�L%U��iF�v[�6��޻qh	P�FɅ�z���H��I�|_WvRc!h�=��U��Q���}	�~6���D�kC�Or�b���Z��i�~��V��+��wTn���e����]>��G����\|8XM��ϻ�d��D BG
9��������,��:^CR�<H����Ӯ#3V��$O��tւ�j��U�Qa����ݏ����U� �V�xF5�J�c��
5��n��4m��cXR�|Q�0�7���R�[7rkͱ8O|���ߔ�0ζ��X?-4X���1�M�"�֗ �t��`/Wwt&F��[�v)���	�>�Uv�͈���Ѵm�������o0O<����r������ڈ<�e���Y�K��K7C��Ұ�r��oM�TAW�]<S� �iZB<����l�{^��p�XtR�Y�?��ʡ��牢����8Єǫ6A���Hs�����ѝ|�D@��R��T¡���od�� ^�_��x��*!Ǭ��+�v�������LK����uer%�Hz��?u��NX�[f9�_\9��m�䙪ֳo�s�NnT{��K���l)�uSZJ�(���׻�	��c/>XEO��4�dS&'
��}6��kF�����OT���5��f��S�FahH��p��YO��g���>v*6�C�[�@��l��'�pQ���B��C��M���1�����2'�خ��t�'���®�q( �Q�HRǏ�(�Ӌ��I �o��pr$��i��$�[��e����!����8��
��[��f|�)�)@(m6���2���S=��q4�f�G]}��	���q�^k�����e�H?ub2;yH~�g!���(��'<Ia�>��X�)un�S���Ac�O��4R,�H��~����/f.Wbs4��{���P��/�����O� a��q�=� ����Z�s�ĲUu�WDJ��ݶ��0#���_J�s��)�'���ZCY(H�>���ߚe�GE�Ђ*a�$j
��8��E(غ���S��n�x��i�z�ꀐ��1�A}^
�Ѭ?�ۯ����^S��xS�<A4����"��B���ѻ���e�3Oǌ��t5��Hڥ;�Sf�U͈�<VK��3#Ӌ���z-r>ו*�^d���5��Z�n�.��[�ő���Q^m��ǀ�E�P��M�&F��CQ	!���,�	V��7
t��sh�JLY�-$��Yx����|�z��K��,̱�>|�2�n�˒�[�y|��n+�å�=�6{�F,��t��G�8���8�Z\2�V�Vƈ��O�5508�T��D�ȋ�3I��H-E�-c
�x8/�	բ4��H��[	��!�'��դ��� {�ehD���8��;"<&����R�y����P�D�1"G����q��Y.׊�7F?�fb���{R9\��}�x�����v
4�-���Q=E$D�e1j �e|�;9���%8j�x���,�9
�;ev�� �mԳ
�a�3�O����Y�1ZLQ�
�hL;z埄]3v4�Dz��"
 � 3bW��DO���lZ��ת#�`�c��y�R��Q��+���M���dC����u�m)����ұf�m4��ݗ:���	]H��:a�ȩ+W�L[����a���49N�~s_�v�c���Z��[�u��/>�y^�Rf�g��V7S��H�e/�T~r����E/��s�o�i:Wƾ�SHZo��Խr��J�ae2�w��s���SP�ß{ԩ����v�O#=�]V�}��(71�O�kb�m:�=c�ۼ�H�ǶغEsﰘֶO��,v�֍7�-�3"B�ɨ~B^^�"Խ�x$�+�b���i�q#S+��P ����� d�˰��;?�ڥ��Zrj�?N�.�q~b�!Mp��\�V����+j��;�9�5�\-0l�c��!]ɩh�&$�g��Ԥ�7Mrl;��.}��3%��=��
 &��-|1�vG����
�K��2�����V�X+ᧄ,?���Lc��U�Z�6w?�.�p��w[�i	��Fc�sfV�j��9��C^��π�j�l"Y������B��.���#-��4V������u��`F�b�*��*�6��a�8د��Z���I������a����u�*R�ƍ�R�(/�i���5z��?`�v���"�2U�����IU��յғ"�cgjЀa���C5{�s��R^vf��Yc�\��.�����(�[H�� �ӵ���F��o�w��@2w��J�1��̤���2Ӕ��H�e{sv�<��Er��>���e@�3%���ǑPˡj�p2���
9�͚�WiA��>Ĵ�4�#��喂1t�Ԟ�<�C���>ҝ��P��U���O�I�c����H�KBa�vOp���T �>8W�c� d�gw>���!C��K�Av�²!���Ȃ�Y����������;I��&���Z��y{o�l�Ջ��<�+�ܷK����	��	Nv��h�Q�@)D�,شWW�v����CQ{�>S>��[l�Bi��p!;�}Et��1���Ką����Q�����3����ks-в`�d�Ȧ�Z>�F����fws�M��.����w�9/._���o�Z�78x1ZX�8]��Bj�\�5vu�'�_�7���ŶyhE��k�����ϸ�e�9`O�ڝ����o	�>��j��DF�3�}�b����WKf�m-��}���͵Z��� .vZz՝'��D�q���O�|�3�x����`�R��?1�T�1�X@o�c�W���ƴ������0s�i�C8��;�� ���#��J����v;�·��E6:,�\G��6x��Ȯ4��E�����D}*���9@���ǓF�e����Y����g#P^�͞�W{8H�^���b|�,�aL9	��UA���ZG�pH��#�y�w7�bU�D}��LFX�T�gk`��L�K	"n��M������p�cc%*�Jn2⒬ʇ15��+W��� �>-P��V}ܛ�� ��i}?ME�����ӛ�vd(1��&� �Zn�N�MW�賕4m�.0�(�E���<j)��b.�&�aTf+��`�t��맋@���d��5��3#.���q�� ��g�Wy<�X���Ch?�`��xc�QJUMǒ��}z�H}��b����M�gm�rB��?��|$a02_~(�ɟ][d��m��.U��KOI>���]�����ҥXJ�������P��0<�bՄ��f�A\�Zg{�f�Q0��:׾�{���C�;���G�媹R�q�s�n������B[��54v�)�뼝*�:��^�~�ZQ��5�$�&���W<R}��U�dC�?��V��oM{-=��9�����¬�Z���| ����`'?�d�*�:d~�xl,Dިi�Pn7���9�Gm8�S;��C$+sҀ�B��`�@d}�%d��zIYyĂ¸?1V��Q�Z%jpPOP��~��i��7�vO�(����k�	.�(;�uIÿ��ʥ�b���ge�b���pD^AK�'�kI"n����'a�B��"=��c��Ȯ=.�h7F5s��P�r[Γ2�A��y���QnaPJ���?��W��}Ҟ�m�%�Qjiq��df��{U��DH��W6��y����5Ŗ�~��������CKܒ�[�k�w
�z���L�\�Fii�k������_�qW�����W��`��� ��eC���5�mY]�����M������� �&J�>5g-�|�(E
9�`+?Q�tu�
���G��1�=���3�1x���rޯ��~�0���%����\�}�y{�'�i ���fgV�!p�ߋ�+J(�;��3��~��/}@��l��L^rD58����zc��}�v��X�\�*�r����T���iy?�	�$V�9z���ػ�jdD[�YY����`�D����vL�F�
z�ǁ�f�:��R�F���!�np$PO{���+��@'����q��M���:���������ʖ��Yi����B�q������Y�K&�LEZ⤃�L���*�%�����QzY� E������?��6����q�%�ɏB*�-�s�թ��KQ�v*[=��O�/Zb��f�/��J�[(��C3��?<'���� ,6:i� �jً���F��i{©���Fs��W!��/l�F�j8H ²�q1&�y�"�k��f ��H�	�Y��TuD�I�5~�z�ĝE*f�P@a�����V�٧�� �\���"b�%\�!�����R���[+�ˆ��ڹ �Bn��cw��I�7����{��t�A`�=r�-R�R���3��XؘV�B��Lz�T���u�������\�SUȜQѸ0Ч�ϫm|8 z=[ی�Ը�]�"ty���4OH����g_\�6v#\��`Ț�c%ow�I���A����zj��������L�Y����g3>�5Y��!�|5"��R���[U+������ŀ��Qr�~U�Z&�3��a�Ak�:#��I�k�*����n���)� U�J�g�>�����^���q3�A�HH�{i�ެ
9�!;�n��S�Jͥ�d�Ř�,�C�k�k�KV;Q��pB�(1L`�� �9�+��|�ː�q�Y���އ�k�� s����=�Q��-�`��T(I[��F	چ(�޹�׾���7�)h9d���E�&����0�L�C�|�������|��@�㄂wrXҨ�;wi�����b�b����28�`�R�&8��-�,����6B��+EZ��a�O�|G.g��dm�j��srFn�1����HP*��aM���O�R��`6�Jk���K� �l�AW�;"b2J���<pT�%�X��Ua�A4@�|Ɯ�G��;�k�g��t�+g>���?;�����Zr\	����Q��n�o�F& @�<��P瓬�wUw	p��u�-7�¬�x�ق֢��p����!�*�����n5�J��@�5A��%p�gW��u���W1���X�/G���#&����.@9�F��!�����ռ�`�� �Z�]커o݄;�ȑ`���c 7v������6Ԣc9f�b�����Rw������i��mJ/.�/���4?F�0�z��D����olO瞌,T�1-K`��R�H%tb��@����2>��8�tmB������Mj�C$��Țn�O���k��Fz4���2��c��{6wX6}��n���X)co�����Gr"�� g�S$���Đ��1�S�<���0z��v����K��o���~��_��v�b�$x�XY�1�����Y�]=hk&�8��99@�w	�Ovz~"��Ak�xoƢr��ҙtG��2|�8�4�[n��7X�rЭ�T����~�CM��� �}n_�Ό����W�� �%|���/ӻ�L��L!d=�u�+D|���xQ�����JN$$����I-�`���]_�
��c[hڐ�w|��q�$�����[�E
�:���}?0[�.��c�Ѩ��"���ɖ�T	=R=���6�����Z�'�?i������]���2�;F#������\�����.|�F��:.9�D��!·<�n*	tY��0���l:]Mݢ�#�0�x~���^���r��o�c"g	�c&z
.W�G7��M\�^���o��}�r�������}�blHߟ� ��y�4n����4�0�raL��Ur������#�Q�^�b�\���
{�P�]����I�U��R����9�.�>)A�Eם����9�ѱ4%m���,F=k���ŀ��|
"�0wߕ�]����o4��wn:�J#�XL��>$�%$�8�I��'?�L�'��J�k��5�!�^�}v�MG2ZX�9}�i��_�G9��Z��ԭ�'�uχm�O��Z;��s����+�m�2�祚���7���k�ZF�����C�t����R��C���!�]��^�.7`5ol�h�C;�0�_���3�(��&Q���βR-�	'(��3����T��"i���GS������V~�g�8u�u���N}c�	�=N�_RJs}"[y{j�P�r��C�����oG�E�{��N�����$b�CLм�B1d������ii���ќ������J�e6N�0�!y&F��Ew�H!�ب�K^�4Q�6�&��H-�6z(�[���4N���밅le��^O��T�(E|4I�&1D��ShЗ��g�I���W�P��F������2�qw�\��Z���}ޅ6:��%A���EܥA¦a������.ʈq�GX��˞��Im�1/ץ��/r��j�m��i?�m0��$!�t��ʁ�w]X/|'��ע_���[-V��w6��/����o��br�,�J$t���s&�o(�J��
���>�����RA@�Ƈ�^���ܧ��d�t�9��?S`��������y6��WZ1�l	}d4��-�!ˏ�2z����z�3)E�<X��}�;Fb7V @RW�{�h��_��bӿ?,����G$����;�w�wV�T�li���e�_�� �����`��3c��[q b��~R����+&l#-��4����+>���l[��B��콦�WFU��8�=;�~΅��O	��6MZQ*�\�G|n�E��������.���'�����^��Eܡ���3�vF��7����{Ý["_����(���u�Ŝr�>�Xk2�ܔ2��dq񶻇Y(J%����j|۶��t��m��d�v�C+�^ٗm�'�?� ��6�a5��˶��>y3�Ie����v+5�Y�?��o�}�� ��Eޮ�1�Ƿ\���O��o�����D���,a�����Ih۩�B��#ţ�_T�AӺ�L�cU����/�\g }��� +c���@(m֐žė7n)A�>����A�od�����B+=��烪U�nC��
�(zZ�$v���L�ˮ��yxG!��Ga���kw�T�u�!
OZLLI{{���P�PB��_q��}�EA�s��d��ʙ�żЕ�5ѥ�sO2{�J��m$P?ބ�$}��	��y+�yu���5�jF����
��X�&H���é�����-��` w�]���&[�}�h ���<T΄��qԊ��9<Ū��lm��@L�A
�8υ�~`Ef��ZsV�_�~��|ԗ.UR4�U��Ƅ=�"B��J��"V~� �+굸"�D��q����L����R��Zh��7�}��I�r�r�l>�U@u�l��@��J�b��yy)և����h�ՆQ��#�Ұ"��7�֝a�rd.���Q�{?/ٓvc��* ��<�Jt�RW��f��]���|'<��/Nx����L���_��0�<��¯��K�\�E�c)O��$G"�`�{K�ZR�<��ۣ�y��d��Y]E�CyH�ڒx��
)5�0�����nU�dy�m�H>�Z�S��N����l�UQ)cA�LhCh�G�>>�}>4CkZ�7�A�(R�,Z�8T� $�IȬ���$=.�#-<1����C������_��&�mk=
������}��vG���ˏ����JĪaeX`o9����j�v|l�V�h��vx���� 1~3\�.�Q{W�b�KMŪ�n�����ʂu;	��?�0b�$�STU-�|,A��r��
4�%e�)��b�P���BPiS!�9�V�w}{4��)�o�Q���1-��?E�m�����2�\�Gg��P��}
���V,f�<fa�=�-�RuG��{�쁂?-`)��Be]^�-:C�a�랕��IU��l�Ea��ʗ��F���Z~�>����B��Y�.Ϳ����r%��L^^) wC����m����Q��#�1v�uC���-�H53���-������N�-��ޙ,y��J&�56��H$WO߆	.fQ�.��LWm,��ݗ�����B�:=���Ь�mx�[��vo@�p����j|k�^��.�VveN���T�sayN�/�ԅ���H!>��]ip�Z ��ʯ0bx��5ZC���.F��{.U'?���Ie�T�\�,��/���s�tځ�оެ�%i՝C6�`pR�&Q�ېryq����M�Ä��,y�Cf�gߖ�+p.v�� g��8_p��0�mr�ic;��
|�^�ƹTȻ�Ub�뫝��up1'DI����˜D�s����^���"�/�&���tW+{��9�%�"�����e���=�a��1J蕕2��{�K`"�?�=1u�Bk9Q������u�S�$���8=���uvE	�E99����w��:3����g'�$����g��S�G����v�Jz���C�k�uo����%����J�J�}_b$d�t0y)oX��ȅ~F�wP���3I��l�H+��>�Bނ�����L�>�}���}��Lg�m�%���/�խ�m�Z�&���:�: �w1J�����9 ]��4�$���n!h-.��H;��C� )���t9���.���3�]�-��7���G�,W�K��0���^M����m7*
�r\a���qe&��wg#2Aq�*0@[b��*���HF�����o���mhk����=�n?Hա���F�R���o�,&%�&�$_�o� ��Ε�f�����,g�*H��u���7�w?S�+���J�?������9��J���(�C�0gw��ïW�>O��2K�p� סē�A��~�lJ�s�M��n�8!��E��9@L���u��r��B��tgs%fm�Al����ӾȐ�7���GY�Of$T�tJť��ḫ�����SM��a"�ȕ�G�ΝJ�@6��蠶�A;|����=nDֹ���]Ŏ�}P;3�J�W��AS<�I�QY����-�DU����`�VF����S
(o}T��D��z�t��� ���Ys�S_$�`�1��wB0�9�'�l:�.?��e�[N��y$�u��o�@~l"���1n�,�3 ���pe����t�p&��9�J���Lc�Rk��b�P߾�4���?���!R[㉳�7�����'�_f�-����(�٣+AaP���ǁ�l����e8dt�����%�"�	=����=�D�:���1�h�(��)�!�<����wu����~el�rK�A�63�U'4�?:���h� =��շ뺲��;!�W�B�es��Y��μ�v�� �.�3lf�F������ϳ���T�^�O�HX�'�_.�1(�~�ow4_>��5�m�����M��wm�_:Bt��0r'2��B~��+�<P�e�j�v��I\ݭ/V0`�۬��Ĭqѥ� ���3�)?��Gvǽػ@5l׷y=���dx��~�,�+gC�m�\[0pU���]�UI`����@e��~*ځSW�C�� 3zzjC  #R��1!�0!������n'�6�|T��f�H��.r/�q��֢U,d�W���4�dv�F���[]'�rN ka�A_l[�qY�;�ՙ���A�s�t ˨'d��ퟎ�5��k�AJ�NϮb	�c�[�T����Γ۳c��! ��xc�(��A-)�F�F=��x��e�����3�!^T��_�=q��C���s��f��I���>��Ϋ���ʾ-�η�ÿ���*�m.����АО��\���'�-��`#E.��|Lg9_�f�U�>鲢gU�>g�o��	w�7��\������i$7��h�ӭ
�9I���u���O6�;�d	J:�C�!�x�m�5P8<�Ҋ�{sc���y���9�x=~sv֗�f<������/so1��ccQ�T���e\&]���b�|���W&"myu��0,�C�q�F|���f-ٝ����.B\N�W�n��fD<59���q��e(y��{���qKS���F�V�Y��$�q?Xceo�ߤ;��9U8��sZ"豴׮e�Z�'d�@��kU��"�[����{�k�-������&���u2ض�*����|-�K���8�[my�dPQ�aN=�3���0�z�������`��"�?���޽�5M�^wmg�ӷ]/�Ȃ�LV�:a:o3�y]����7��b�������[�]��'�����Y����w���-�|8./����8��Z��ϧ~|�\^��p�X��;�a���x�{g��'�	�^3K�hMط,�5/(���c"r@��Lp��;�c�r����&X��,�Ŕ��YFp��iI�;6l�[R1�L�A�)����dA�0�����]�dt1���;�oݨ�X��.�/�p���>���THK:�Sntm�"&*���d�@L2���>)5���SQ����� F�/B����P*�ޱ��HN��_�Z*Y�<s�k��!�"N���H�	�=e����naH-t�X>t(t
�j�M�A��߻p��,�F�%-ٗ����(��8{��I������I��D/ sn�E
ۣ��]7�n�n�q�'.1�7���?+����M�f%z�&M�9��U���aű$ht�|�k���/bB��zI�K�v��T�G����?������8ߘ\�<�y�Wx]P=��1���?��^t8Ȃ],(��&BH�3wǯM�Ǎ�>���:s��%�Yk*l�3D6^�!����45��v��	����1h�Ɋ69�TɑaD�,deL� �D���7���Ȗ��@�����:mL��<v~";�����-$�ce�i��RK���'O�-���[��-JX�%���U��x{G߽���&1�������`**� ��;]�&m|X
�e2>\�r�[[����W?�\�]&�T�?ą ��q͝{����2nk�Bu�.Fo�O�B(3��J�D�U�I
\!$�׋�/�ް��'=��t������G]��WP���m�H��
=��ж�Z7�����h��%�C
�?R�5'��!O�/���[�س�?cѨ�H�� �o��Ӫ�D���Q�-P!���e
�[b���-w���*��>��v��#�OrȌ�9gp��}��|'�!���� q���������\�w�Z���;#�MFl����}*`��BK��"�O��ΰٙ�ajZu��f M�n������ǵ��V�o`7�hX��)�L'4j�k��h��)k���xc��~�V�"k�����U���oH��-��r��!��A��<�P�'E���+�������i'��z��m}��7)�t�J�Yӫ�W)��ǀ
��񊴐�E%�\�4c��`F�����S�yUL`-����?ճ]��C"<Rd���,��4�I�L���ɲ������1�}noL�&'��Ok%���YAZ^�2��u�Ҹ����g/���7����Khr�v��oʙ��`�YK���))���a�/Ai���y$������rv�迥X�vW����b;]��}���|ޏ�..LCF
�`�;B>�Г���%������9�X3%�'�����BjȎc�m�WlP����xe�JV�l��߇�z��.2��TW>a��a�2i.$:'���e��rh'-�����;��A��~>��R��[���)�#����J��d���z�>)�\6�45�|��",�d��8�2d�{����4cNk:�*�{�u��p��A�볥�O!}a�`�/\T�h���K�V7���&@G�妋07U�!�$G�Ä����q�Zo�#���
a�\C���n�*������5
I}�^>C��|�֭�a*&~��-Z�nL�L-�� lt�ߣ6&ϸB�+r���XL�������w����cGL�Bz�j�,MI0/��4WW;���O����FK�$�Q7A�%E���r@�+Ԓ~[�k�jF��IB�`�+˰k��V0-<�g�g�+Ի� ��w�*d)n��=ZQ�']|LL/Ip��7��>�6@������=�s�a���,7�@����RH�e�t�S2���ef�+?ܟk��AK���"�n�O�5k����������*m�)[�����'Ϫ{�g�I�*a0��E�̊4�W��j��ހ.F���{\u��@��Xm� ���Br�P�C�.�x�~�$�#^M������U�K��`bj�m�ް]<�]�.=�Hٶ�X��h���5�#�4(��vO$t�y��Q�"�B�TQS����?��ZO��Y����$5��O7���č��N^2�S~��������B+D2�����D{����w��WA;��%q�l�}}q?�hG���usb��.���P�x�^�M����xR:y�@������'���+�{�#g�:�(�ř2��'h�a�/E�;�����Z�JB�p�x+9H�6��`���� �}~�����8�3��N�r��i�%��I��B׿_l��!t�Kz��S)�9/���źN3���W��p���x��_���R���x]����%'�)��b�S�.�W�y�T��!?FL�1�`w=�J��p���i����z����O����bX�S�u�\�`z$�a�b��C5�K�����[F�,]Ã�������=hpw$XpN Xpww����������?�:����v��]=m��R���nI��/�d$���PǞ��6� b�덜�*Ib���(�v�����*'C��B��Z�1��R%?��J�ǀ�� �Ϛ���𦶠�����ޯ1�8�J����G#���k��4�[���n	\�e-ЭE�#yZ+.��̞Z#,���@R �#v\D��� �	�3�Vm���R>c����H��l��on�J�'���[#�y�A�ᢄ�2{3�
!y�P���G�LĈJ��}ʔ��Q`��Q?|�������.|�oɔ��߹�mr�2��zlT.$��`�������;c��3��W�#�:����-#�	^�@d;�'_����Tt�[���ۥ7z�%QS0�J֛k:f�N�s��v�^��#�%���?1�m���d�fO�;�p�f�d�p��fZ�FS�AܱcЌ�>E����r �j��M5��gc#��%��wzٝQ��l�k�u�m����3�ɸ��3_<�v������l	��st�wS�+̏�V�f_��M���1圜�%�ٛ���o�\�tnt��R<z����W1��w�e8�:H.���*Xs�{������fw=�>�[�k��u�'�E��J�4�1��t�8�S0�G`�=�x����nہ�k:�Fa8�	-b��g��W���	d5E��=� B�T<v6>SV��������$���8O�8{/*����$Fd�h�f����Y���ꝫ��D��6M������x~��k�%���F���_]��d�+��5�o]D�I��B�R�6�<��u>~�T�����Y���-f���Oe�M��2�Y����#~|_v�}�+e�-s�UN�C��A �鈌�D;nN�����j6���� QWCJ���n��E�ߙ�59�}��]�힜�_�������0�۴nf���L*��I��ſ��!y�W˪�b]���w"��S�ؗ��������o'g�`s<���N��l�qb�eҊ��#�W���K.R�דy�gdy~����؛���H�C7@.���o
JJt��bN�[b�?�	s� #/��]�p���gW�x/�`tFy꼝����������'cVc��~�Ww�f�U[A(�V� g!�\��ʹ`��-����]�Nכy	�����U9�`�4���s������[�w6L��������vX�&|��Q�΀���՚�b5�lJ6��˶������(��N��19�n���?F���ӿ\�/0	��h��U�m^O�CA�XJ/]NP4�,'^Կ���U2�͆�Y�B����g�y�<�K1���|Ϫ��/�rM��q_P-�����C��"l��`���U�p<�"� ����R�ۛ'&&�OoG֌�E�S ���_���qZ@�~`Ǉ��I��P��r�~����2����]NM�A�m��z�+1`'������G\�G\�k�:�~3���S[g�;(xrZ��y�z�z�ƗR��xee�b�v�1L.�%� ��Pu��]���SK�AH
�3)''ʁ3ҙ���L���[��~��|m��`i��kZ?�oe�����{1��:K��5NL�Y������^���]��:�9���S�g�y|t��F�1�%l~'d�$d� l� vBxǣm�MH.0>"��l�G?}�t3C��-tc�ﾧy��1�k=�ն�WE��u1o�����~`lw����:O��)fm���3'OȠ�j)l�!��z�gd�����)Q�R�绗��`-/�'|�SW�O���;]�}-Cl�.��f���������5.���F�L+γ�1�AF�B5������/�릫U5#���hI*-�����5�;�b��E��A֬����=�-�S�*T�޴0D9G~a7G�B@�um��v��� O�8���ٗ�"�#�AZ�!��w�e���5�"�F��5#�VP{�z��qoQ�.�+��t����]#Ԅ\>��x9�[K�S�G-��-3Y�W>�7��|���0�Z{��F��6V6�#�pn/�|�W+��?ؽ�M��ћ�u5��h����&���ր�8~]�Q�ύs���#�(��|�R����l�e���5�'nB}�{�\��!9t)~T�]�����)�����TW_�u�h|my"lns�E���,��S� b���2��(jvD#�������o��׊��^Y�!�<ҒO�Ee������#��l-�mh�or��9��������s��h�%�Nc�L�}�Ȏ�f,"vy�hjR�`�N�0=�dLV�)^�t��3"~�c���:Ä�� e�d>�vV4ߋ��Wȱ��Wn'��/��UcH;���g�B4���͛b<%�����@���h��2�A��_P`oV7A�����i��*#)��g�N�o9�ʣaT1sEOy�M�u���Atoe���jħ�vX|���U����X^���]�m1���$����A�.T��ԙ�'���� �K*�\ĵe,Pd,@'+2��S�k��F|Sr���C>�9�W$"�WRBu��L��	�g�A��_�, �B���Q�kx
׍�߯�ս\J��:��[4=��U�j�`@i8M�����^�D;!	
��}xO�o�Aپ�-���u
#ᳱaI�ʓ��!m�x�֫MA�QS�dQ'���ʴ��2��69�P~�cU\#!؟x��ۮz(�)��F��kӽ�o�߫��ik�D�dS=ї�
�m%��&=u���PL�Ծ�521YY+{�������-6"��O#�GG�����/�LmYɌ��� �E�Mx՞��f�-�)�|ĳ�;���"�w�R��t��W4qH�.��8 �l^^?��������͓$3h��_�i�Ah$9����%N���%8��d�Uّ���AD��*۟?"�YW��UIF�Dj1%%\�%cd��9R��N���o���;��Y4��7׿˰8Yаd(�� ��o{�
������.��e�@���Ō5'�hJ���d�im]���Sag��kZ�^A�33VSQ�e�)d�f��=��(&��L�<z�2�Aj?Z$�+��$S�dlѻ�N�K�|qHy	�w�/q����1´z^��q���d�O���(ؗS���B�������,e/H�P�}H�I��<�^�)��A�{V��>@^/��T��� �w�E����ܣ�Kz���XV(��}�؅8�cLv�M.����2��F���G��,.�[t��bcK-���h�ⴔMe����d��O�e_4{I���?���l�ުW͙���u �F�6�I��ǌ��m�!���=t�`%��\zԳ�FBm�lz�Ln�S�.�U��ԕ[*�_�#P5��S����U�TX�%�[��~�㣟r�;*Q�.�h��ݒ�i	`��F\ &�߇:�Pء�>"@Θ�d4ЀZ�t����gg�as��E�,m���?�>�*��3�j�{.�u�ph,1f6����R�'�s���d@�h�'Jp��ښ�*����@,�N5,V�	~��`(��O��Z�m��QK��L��j�KĒ���X�r��oV{=��ֆJ���W�2 �ўa:A��o}20E~ak�Vᴍ��Z�Ҳ0��d�S@�\��J����q�&&n�U���*Dl:��K�t���`�\�E�wE�r���WB}rɡO6���������6s��g,�ԙK�@��&Y^a̼2���޽�Z�*f�~��u6���i��ԧf�|$��t܉;����2;���?H O
�@Њ�y�M�GP�6ӔJ/c�}`��,)B�I���i�݆` C���E���A� U+.�ʕx���ҧ�˕so���d3�=��H���g�@�cX�lN�L�|�n!�L.��>��?o	��o.�R��@���$����/^@/�Q��˰P3��k�T��?�ǹ�Ͷ
��rI*�GK��������J8p�P��[3D|�������y���/_˒�Q��T�L��Zr�O[(_X�Ͻ�h�^�e3��4��8L]"݀i7��!���‼�¿������Xܿ��!��O�w	T;{�M&-�bt�8��7]�ʭ��	���Q�~�!�b��b>�s��&=3��{�T�����+KsܲZ=jL%�D4-��X@���[+t׾N���in�"C&t�Ǹ�^w�]f�����e_��:(*w����6O�P�e9�7�����+��L��b�(�mĖ�����?Ι�I��������x�vlff0ϔ�TZ0�S���>����Ң鿫hݺ��#m�Akhߨ��흽��
o�wϗ�Y����%׉U�T�V��|Ig}�8v&�|��L�q��U���3���5�W��m�-p���n�ħ1�W�;6��,X)���LE$(8�!�2�-���VP�H����F���o,��e�Vi������T(�l�ڨ��3��l���?�4�ٞ����F'+ʶz!�}�ne5l�ס��z�Ұ���y����n��eW���{�{΢���)r��.�uQ���!;߷S�i�`�B�l:�d�S_�m.T�:ۏ��8�7;��e<��b)�kp��D��:�Һ=�H[�{H��RU�N����~�Z~=��-0�?�s�z���Vc��M�ϗs�U��/����L�9Ev��~CP�X��n)d�j�>M�
��U�q2L���� �=�3~�W�C��s����M��ҶH����6����J��L��魗�^�ˏ��|�򑢚s���,���~���Fa9t,�|D�=��8/3ª9w�.kxT�[c������a8ѽ�Û�ն;׍ԛU�����J7I�c�sJ����ޓk����z )��$>�|B��¼�ȶL�N�Y[��z�f���.��c�yH!:Ņ^>�t2�DOrO�	1���!u�����j�#��Q���%X&>{^=&>�(�֠��b�?�Y��e�{)'�:�5p��[+�)ƿķ^=��Ԩ��~Y�B��wЃ�c��zk)8�7CjT��ኴ4��Q�����PZs��ع��Y�5��������u���*�'�r����k�;�ƺ�^��b��]�K~�_�xH<��=�K��B�H����K������y�o�RY��|_8��
&D_�6�6n �/��_u�徣É��i��l܉oڿ�NL�p"��\�q��׮|�������۫5��'�Z��I���`�{B[��Ids`BTf��& �|a��Vz5!��jdJ����~zE���DZY�i��0�fT�NK{���bo �"Y��	�����3�r|Oߞ�F���ڷiB]�P����K�݂�s�~S�+w�e�Y!M��o`�U�_;.��t0�n��n��{<n�~�����OY��J�=�0��� �����������}e��E;�d̈�:�b
��gÕ���plJ)�N�����ߝ�_\�8�����2v���c韧�52�rӝ�o����|����	�u���B���/�=��
�@ �X�mS���R�f!sy�A%��M�ѫ �"�L4ǑԴ��Mc��3�������WRls�'KY -Oy�Y�i3�i?�~Ww�qB��1E�*(G�g̛�n�+�����z|�6!ľx_���{�π�s��0�wߖ���$���ɋbOX-��Z��S�v�]�w�Uc~�ډ�b�O����v��V[���7=�z8��:���b��
�1��ʥ�3���Y�Ғ{y�tUo_S�=�^��x�Rܓ�E��V���t��[(
f�� b�*��l�z���b���'Լ������ ���<djG*�$t��*�u�kr�����g d�� ���u!�l֨

]�L&>-Okχ'_�T7.����z�h�������o	X@�J��"Tg)/x&S���Ĕ���QN�θ?�K� )��}��k��-��Ѳ���&(ǉG��p'$H���3��:��_�U�/�$�E�(�������Sz\�G��O?ɷ^&t���|
w��%ū�W8s>�/�];��8n"q�ޤ���&�qh"A�6����DT�X;;�e"B�8_%-h�s'��ʏ	��É����c����H�d��s����^�&I�ѹ]ٝ�����e�-[m�q�M����-�
�����:tR��J�-O{9{�ө��.?�V�ϸ����'Q�q�����Ɋ{=y�^k�r�$}j%��A����ű��e-ؽh�i��y�|�qq��jY��H �۲x
6���ò��7�����J9X�����rȩVQ�GMX+�F�m'�5)���d �%/%d!G�z����ix��j7+P�E���Q47{��H�=	��B�N�ʗo����V�R���!�.鏤]B���<Z�̙)��g'ށ�e���b_.�)� ���~��[�xEשz���jӤ���}n�S��'�D���������*#��~ik�*He����e�Q\$m~��CzB���W*��ڗ�����kq���m\�ɳ�P��OQ�����|Q	Ũ��᫘:�n�4��i�i<�>�S���+�u�z�?y�>R���ԥ3�k�J���+<Z"��x�i�I�E2ђ���s�#L�Ղ0�˿�v�ޮ��}���+�����1��_�M���@{�B6:;w8�M��=ݻBtZA�J�r%T���J����`���Y �N� \�_�+=B�|:p�%<<��������E1�#n�2����p�v�;��P7������K�*H�i.�#簈:�ބQN��=}�*��hl'�r���S�����\�p��-���)+�q�ϛw��~?�ヱ&`-U �P����@5�/i56���qӫ���ul>@��V�RzR��R}����C�`@����� YP�#2�@w�*̅��3",r�W���ApϷ`G��f����X+u���|����U�c>�1�N����Y���(U��t����/��^r���J��\����9(�)�����vFif�L.��3�Qy�02���<���җH뮞<RIK=���֕�/)�4~��֪(���§��
�К�%y,�&���9��qP#���%����1�Y�t�V2�K�:�������0��Vyx��������e/Eڈ�1s�۳]A�J��	e�ķ˞�<ᴌt������`P��k�z��WU8�&���`v��7�T��@��Ć���k2��2�̏�w�WgQW�*��$�o#����]K ����[J�L�'ec�t~6��פ��JFDN�S����6r��u�M���)4}�dU�MMZs��4&�<-�y�jB�m���3L����c��H�PQ6}\|�r����E�Ŭ-Z���p�t�k�&�[5}��5��}�8`w���y�5�����&�`c�A�Ʊ7��Py?R������2%�:�/.d�Hd.2�s�_�=��76�5x�B�_���Ra�MN�iR��6����~ٯ:��,k�𽇃M�.�FNG�O�c4�+�($� ��Q�����|]~�9�WHh~~m�Q�;Fi�P		o�ҺX�C�;c�r�p�u@���>�}�z��h��Q	J'5ux"
�w1%qsa�?��ް�G��吘�ż�����lW��5��&����-Po��/��(P#b�����f�--e��ы��#�d4?�ֽD{T��Gr�s�^^)&���)���iQ�Ҽ�[�.�>��ʈd�v~��#n𩭻gzo���$5|���Ԁ�E!8/�n�qhs�]t����t����gc`�����Z��H�1:��˒���>�z�4횊p����Bf�zn���	���v��	��HF0^��^! �R` ���y������*�j�Mh{a�𩖧�8\��dlO������!}i���WG�]-Rw����~�����\�|j��a�O���>	�.g�Ռ1�����i�?�%7c�MzZU�o�6�e%0q��f^�����M�~�Wg�
\	؝���%��o��z���Ⱥ���g_����s7慆��5<��?�bz�������St���G��*���L`ڴ�Kce��O��V�d����.KYi��	�O���z��cߙ��5��OI* ��s�i���B'�(N;K���Io�\ek��T.YlPD�uM0��Q:z<&c���*�(�Ď�,b��1`���3@mQr�`���������~���5>A��B�d��\V��:�y%�r<��Ɉ
~>���Sh%C�jr�9K,�a������5i8�]zvs,1��\��z�B� �}L�P6H����*�/\�ŷ��;t1W�n�|-�Y�֦ԙ��j���ޕ�h�wx���8�f�$�0V��L���#�8Y�����IA0�L�\���c�3_�f�6����"�����C������y;R��	�4��0�H[A����CW�f����>��Co?\���E��Ĵ�7g
p�id��u\"`�@OTT4�;��B��/�Lu�h[|�$56)���ت���,�E�@������A�;b���G�9[�rd�I:��f�{��3����۪ ���X�֫:���:ƪ}:�����%)��;����Uwp��NDn��e�x b�&�o�p
r�J8^�s�Еe�g���8�&� �-����l��X�ҍ~:�3���BQU8�5·@cV	"�I�)�
1#�Cb,m��T	]�٭�g���}��z�ɲ�v�����*������䒷TO�{�y\_L��_�HE���Ay�]d����K����;���_%0z�*?Y�
t�9w]ꗃ��T�(N�慿���U5��%:�"�����cE��v��[��O��*�\���A@�Qܼ�t��?c<�?�Z!"���Ϡ@�T ��8Y�D�l�4���l��eQ��(8d�^��Cu0���7��2���u|��}A}ը�1�ر���fH��Q�ǼԬ��m$��N��7����wǋ�}~-�!!�'E�[$Q����\TcI�$F��c.�@����q�u9��L�G��C@i�՟� ���l+�����Z�v$.?c9"$)�Fe]���_=�Yi�V��g%|�+�As�UR�y�t�/����fW��=.j��kV�v���4��g��yc����H�X�Z�c�MbEg:^Z��t@��'"������l�����Tgw�!VS�����hW(#5�dBa	4 s�h��KO��n(��vL1��蠏��@+L2Ԫ�+!(�B�!EV�a�X���N���੐D�����;���G��w
~�6��+꠆P�Jܛ�ȋz�����W5�.Jġ���cJ2�!C,�,[?tG����fW�{ɐ3�{��xI�y���+����׈�޵,>�$���@c^�M[������)6	6�@��ܥ�����x"`��m���M�5�m$��͛u���8��� ����W�j�z
���v�~U~� ,nN8P Ԅ�]3���h�J�����6���,ץj�x��n&�	��;���� 	j�ٜB�� �V,�$l�G�<B�qܽ�Оj�[��M/��!C@��	𱧁]�_�Y|�3��r�k-�!�]�̤g�~�ط-g���--x�dR�u�e�2{�P��Ix�C돒���d�;uʌϛ�ס��'��{�F�������a�$(����'�"F��Y�0	Wc�:�8.G��*�C������&�1x�p��4\��lbP!�G�c''�]��c=J��Ve�4�蠗�5M֕���p�6T�ax]�B�s��IL{��d|�󃆉�-���#��[JA�(�>�g}��CM��� hS0:����[lpk<�{��Ƹ��A�mbJe��`/���UT�\+mC���9��S�'���e�������<�����f�)_��[�e\VUM���r%8����K�s{�L
	�I<?��J���^�{.2q�'��M�.��, L
ڝ��E�T\Ο�qqhFI��@1]m�*郲�/��|�?�7�I��f�T�p����E����C�P��3���Ԉ�rb���6�S���<ǁ4|�P�:���HJ�$D�S���?H!ㄱ���WN&��#�x®����{]�b�G��h�D�hZ�tY0.�ew	�G����h5D���c_+IqR�t��TM����ϲ��(�[ը�}'�����}���C�ɉ?�"���a�u�%-xu3�J���>�͖[��z@�Ȧp4�b�'�vQ���z�����ȫ]OI�����r{���x(������M|��p�ts��f�LE��D%ASj��ĉ�-��xm@[�WṭjXC�%j�\93��Q�	O�i�.� ��|���KO��?؀V��n��S��kz�Q-��JǴ�g�����sM�ͽ��2T%�'��%V�-6v,G�(�:�$�l����:�25Я���V���ڌ	�>�%�	'��h)|>{�N�M
�ّ���P��l��&h�Z��Z~�}o���C���b#��.��Y�o{�7m3�9��37<������y��R�ԟ���s�74�UUd���E��r9���?��n`U��L�)E5OS=�_�(�o�b�r��hn})�����F��A����B�R:p3r��{��v�����g�W�t�c3}"=�WgB3}v�?����l������܆dY� D�%4������B�H�x��%Rs����8�>�NXmU9��ן/��tT��ƒ��>��I]�cC�ӈ� �ƚ�U-g�=4O�m��hN��pj�s☠��i�k��r���%N�Y�|y[�7�kD�
?&$7	�r���;���$foq�h��d��↭(���/��@%Ө��^
�勒�����aJ4R��4��=�_����w;����)���Rb0���z�}�8�y��]�3�E���Ýlt;�ʄH��4�I���J��n��l���~%X@k�ꏷ(
3	5&�_r�aU	���EA�U�_c��H��߸ID۬|��$�a}�
/&�([|5ъ�T;�^%������o���e�U�x�h�����Opg��m��w����=wzK�f���מ�;&���3T'���h��o�=�>���'z�@Opn�Z�yU0����n�E��Ix�w�k4%��&���|��}�n�%z�U��6l J.۶h��'�}m�,��=���G��c�{M-DE�%}�L��!O;0p��(�(��!S�<�̋�$��|i������(�`R4�r��	k�7��η%H���7��y�K���I�\�����xm'�I�u�si�M�QB�m��rg-Y(t����r�s5sBE�ge׸ǨJ����Lfq)y�B��Ot��u�6O%`,=�ׁ��EP�dqԁ�»�r�t�u;��1����d��b�/'������S�h4-����|�[�^��	75�0XO�x<� ��<�g�D�>5�[O���G��p�j�:���?��7�����u=�e���@���IF%�a��"�,b��9�b4���;o�����}^ŀ�av�ߔ��G8�?�7�b�y�	�+�oB�Cĵ�}Y�i�?Sbv�#+:�P��r���t� 2GG�����N�c��CWU:�g?u�8�#"�>���=Nl��K�$����sb��b�e'��
�9����2ji1�q�'�\3������'�M���i�О``��Ɠc]�}�@��cL��U�3��<
�2��c�����9�z���%,�R��_a��2c��kkf�S�}�Z��pm
QV-O��MQ����9��/���|\5ILֵ����çN+K�x�_�sɫ�R�<�s�X���k�&�S:i'��܉��;bObNl�&į��-��Ʉ�*j\V5�i6�"�����<l��Ծy�gAI6��T�]��^����/,���k�[A�r����9&�����}��o1��D���C>"�키Iv���.7ԶM���x�8a��Y��}`>&��?�;NMi�q�4��[�B5���ߒ����B���4S�Fz��#������0M�N�l�[/{�(�g��O"�8Ԟ����2C6ʫA�����q�ۯ�KaO��v�ק�#*'øXE�X���X���������:��Q�Z���������v�HJ�\��o�K*�ej�ncu
r����ˌ[��U[�i�N �R?&%�����DAAD86F��P�,g��G:�\Xn!Rɰ�*�"O#kq�;��E��>]�w����+��,m�P�tG��)T62�)ahSb=l/~C﹗L�#<�G�>Z���/01]X�ͤyB_�y�f��`J�\�x��p1�O�Ard�'��2��_�k8n�W�����6V�"L��BǇ������y.�ʋp��ݰ��|�
(�|��Ib%JV�~�ܻ�t���EM��|��lφ'��:ػלg��$l�"l�)B�&B�G�^I�LI��c �.��
�a��)�n�	��E��$�@��GU���铫 c: @!S�x�� �&�����d���@q!�����Ju
<UA�5�Cl�(����I���hȆ)��~	�
-���@-f��s���G�#�V('�O)Y�?��?�_٫^�U��:�_���P@IT<�C�Z���vp���+! U�זvP���Ό�t�ދuN���L`�w^o��Xxz������VPLD����X[���24�?�z�O.���{B»ſ㟑����AcPԻA45BA���`�x����Ո*^���]�9���.�Y/'��f,QnT%�e���k�\�����w//�$m���_��P���)�}t�l�1yx�i<�~��W��)��\o���<w{�3;� A��OosY3�TB0&O��{B*6�o����($Ԝ�r+ ��,�O�!�>\%�H����������ɘő��c�@�ޛ|3��x$�s�����}��I?0v���t��*>�rT7�A�d{��
���=<h�B�q�(^�fGz�W>��^�� Ӗ�U��p�����������
t h��9�Y��R2��2b�\I�K�HH�*I�ƚ!�g��JZh轾��@9��%$� �$��1�Fw�F�!��n� �\�X2���;8�S�����(�c�F�Yԟ#ɱ��=������6hF�i,�����Nޚ/��R��s��� �:��*����dн����h�t�d�47��_=:�aUqC�k�X�k���c"3��vP� ���y�,�f
c�4�.�	&h`s��0�����Ȅx`�@�3x{���aEM�T��A#�ؔx8�&!�\�U����i�<����"R���y�04�"��P��Լ�rj����|-��K��`�AN=	J��
R*��xfk��P�|u��^p���E"#7#��qt�G�j�4jMZ8=Bh���e����]ӧ�d�t���@����f4��[���3)�)%�m�W�)������Z�m��SY���J!-,j�j0�{��!,^y��(%��Mh���t����W��l-��M�t"{��a�
G^Md|Sv��y��F�t$�$ªؓ��O߉/o��T�Im���߹����7a�y_x�	�
�`�[vG3�C�6����	`^�����o�?�A ���/[K{�m���;q$�)~F��7�l��R���p��r��e�Z�m,!T��{nѾ�_�9��E�3#_��5a����KЭ��\�������Q��e��(yd��z��m{�q9����Ø���4琔?�p��F�Өc�IF�)2M�M�u�f�Γ$���8�V�Ӗ)`� �/]�|P����*�Nx�Q��܇f �m�1�Q�{d^�VK¥���N=�d�aNF�^�1�\�ܴ4}�t���S-��D��$�OA�G#��5���{`҇���'P-�1ϰ~��g�`:,�}��� ��/�M�.��VԼ�I��'��J����=1C�;���%h�f��m�P�*���	�@}.�6��&�-��b���ɑ����z��tp�a���d9섳�$���
�h
���"�讽��a�mZq��(��ň �)[.�X=9p-Th]���E%���J~_n�VVs�7B�KU������錞��� ���o<��l�m@F�J�M���_��}q
�y���W��g�1�}�Lb��/���\W���No�}���m��eq���!�$�1��!��s������o߅�nC�L/��,ω��>�>���v��=�oÄ���p.��>ȕ�(G~ ��C�\�BF>G�:�;(N�,̋tۑ�vz:�hmZ�#��}����X!(y)���{��$���`2�`g�g���-u��lh�i��9d	�Ӫr��|q��݊���gS��(��عq��V���>�v�Y���<�ޢ��8'�"�X���2�o�Eͤ��wJ�%6��GV�烦Э]o~���o���������CcL�pN�a�ݒ�7F�p�c@��:B���V7N���+�>�ݟ0���f�L�	l�_-��k���f�?Y���雞�h�\�G�(�q*��{�Z��*���JH�g�p81�p�F>���¸L0+�߅m��p���� �֮��<NB*	B�"!�NA��6����E<^7�:0�h�o0��y��a�ʉ�Į:���UmT�m>�Q|s�c>��n��1e-�����gf��t�˷��5t4��ު\e����Ɔ|���#.w�Z���x�����&| �J:���b�|������n���6Yt��;�2$i)5�Q����"Թ�a7�/(移��r��b���L����8P���:�t�6m�d��7׽c$�`SA=i����>�e��>{ �D�0
:���z�MG���#��1��uy�,�e�2���6�. ���Od��=�<�)Yҕ�^prhm7Q�m���|��)^�I���\&��S��c+��@��,�-+��#��\�)s���pvo5�~>!�ݭH�(8l��#�z���!qɧ_�{�w���-�>��S�>! ��W@k���s-)���f��?�̧m�!�E��"�xY�&�T{(�T��5��(�0�k�Ow��ΆPo1V�����e���^���b ��+����~�R�wuXY:�>df����;I	��t�	�D�h�`�X9P.�̞2E�3���"�������$ c	��ٵ\�>3մPK��#����]�.�nX��B����jN���R0KY��|P�!������q��O�ioB>�t�lX+�Pw��q~�=��Qz�E?NV{��L�x`x8Nϡ3ў�<ॶ�e?0�q�f�i��F_�A �i�9�(��?�y�11&"��ڂx9w�mC�+ɻ��
 ������o����� ��H��A����p��z�K��������:�24u��a�P^	�Om�`�&W�h'�!��O�y `��3��=�	����Y+b����i�a�X��t>��~�, rV�8�\{d�9����;ٵ,#���Cn�v��vv��\�E;�Ч1�׫K<�_WԱ ��C�	z����6��s� p�/+�-�J��!O���`M�����E����M4ӞCl�Y���kL���+�._��m֡����:��;n��2�5T��n^./=�y��ƾ�/�_��0�*�s����D
�4&Q��{��ϙNçv�>v�֩_��F�����O;����md��?qq[�C������Jz·���@��v�y|��0~L�y��>�|����3�!��>�<}�c����wL���V���Jr�0���Ryg��51�,r`lwX�RS�S�= ͙m�E6{TH�w�6�1Li�+�Y��4S��V%Gt�bu^yi{X@�A�
]h�%x���������)�ė(�x/h�w��������!�َcu��7��M��\x��|L�*&�����9�l^���؟���R�k�t[c�<�e� 28��}��~�׈�O?���43X^C��<1�����[]�RPP�ٮ�ڄ��Eb���*2$���bp�� �_���Zcu�2�Ͳ�r�`^n~O��`+%�b�1�0V�̈!�GK%o[�DA�\�������7��>�'S�Bs��3a����ʺ<QQZ��&��	�L�Hť��� 7\ʽn���jU5���Ei�|)w��E���ۯ�[)a$Or�	.�UI�����}��\�po?i��^�`�X�DT�"͌7��;��=ئ$g���/Hd)�B_�{<����ӕ���ʗ�7�8��G�1	x�7� g����f/(�*H�~���b��U`����g�}%h�R^k��2(;f�ݪ����#�43�T�R���hܟ��W5`��
gmK�5A�B�n�'��m�D��;�x6=qj�#���
|L&�؟[Q��ُ06^���N���!Ex>癁�k`z�((��L��'E���̹�ēȦz*���fWGM=��i��$�*�ST�)�bڐ��G�:����m�����;Gd�<ܭU:�WED?�N�wu[�d*uP��%���_!�lq0B���RR�f��Xo�H���� ��y����}qwwww�]����	��!��Bp.�'���w���W�UKQ5�5��}����M0r棽w����<� ^��9���t�>��m�����(P
;	��M �CI�V�|���s��[��	7��a�����װ�U~�T�ꋱi�
1�$�A|v����D�z��u��<�	�\�&ĹfՉ�<�g�'�i�{h!���s�`̮������f3~��w��v���I0;qz�.o{)}ޣ�;)����M��J;*dŞ���{���;�Y�:07X�����n0�N/���[]:��+��E#���D 	O���d�g9R��P�pxY�O�K
)x��F��1(l͊5����3���V2
�
��r��S�G�=I7�\ A���Z�3��ΊR�C�0��vz��H��+損�AO�kjfGUɉ���1�����ߣ����u��a��l��֐�N��Mt?���(��̪��y��\K�O�{�7��[@�I������݀�Aw�1�pWa�8�]�b�i;O؏y�ʸ�o���.� ZUj�����Tt`q/�o��޴�$R��l(G2|�~kg����aw��+�����aKρ��ܩ��33�_�G�@��Z�1���8S���	��p3�W�#Q����TDWv�iz����Z�;~*�}`��rQ�} U�wݘz:������hq�ِ�(�
�5��A ��
>�����!��',`J�r�J�)?r��Ĳ�#��0�+9+r`��Wo�{��CYߑ|[�Ml۱���<2��+]�����*v�`a�d�T������]�:T4��*�+Ԅql��VHɯ�9	�'��NYWqމa��D_�(>n��i=�IJ2b��$ڂx�sHU4��	���=����u1���"%�φIp�ת�<��nrY�'��t�m긯�x�b��0ط;����fS��=��~/��̅7��p����DD�ͩ�3�Zd��Ţ\�`Bx�����}RE��k䶺i=���e}�q��ek����=�V-/m� �'p�EƠI��?dm�jTl�� OnaU 0Xj�f��QQ`=9��c�vs,©Lչ���������
z��xJ�J��9���	 �Ѱ��A�o�򸑫�@��I�1�I��=������>�DL���v��^�&ʣB�tJR}??��$vр�q[�d���� yhhs����Qh1J��`0oX�)k�qK���Y����� �8!�,��.�8j�u0��V�fvW��S�T �EÀ�ы�ͭ�YB<���*p^�_At0��Aex�I�|�^��V������Qg'l�%�/L�w��w��V��D׾��ť�R7w7�Ad�����%,��d�Ӻ#	��o m�˭���M7��	.��q֖�l!&rZ�6s�`���Ћ[�4����a&@}t���mZ�iʧ�o�1���*�g�~' �]���tj\����xc�~���2?�������<��j]	�t��6��u$vsC{��Rc��q���z��zw�,,���_��֗4m"��#�j���5����@>�����ʟ�x�_G�(� 8�ļ�лG]�b(�P0�a���1��ܾ �J�( 3�|#��_���t~�<Z]�A��7�^������b(�6zngf��u���h>�t��~�W�(L)�0
ٵXWU���T�+�㰛 �]�fӥ(��1�3L�������D��[ޔ�P.�!���aLά�֜?�+s�1@��ymm����-Е^�)���'l�)���d���qh�Úx=85���XJ�Ӡ�7�fP���5 #����>/S���vm�?���{�ht����4
 qݬ\*�g"Ш�)�F�*3�EF�ta��� i�	?6�C� ~O�~*�B����C���w���/��H��JG+*[����9��H�S�af�&f&��'���9wKt��@�I^r�U� v d�?J�Xe�JqQFț�Y���Щ���zHmGQB��w�ܨR��u�;nЇ�qh���a�\�T��˅�������^+l�N�,7è�������e}�A}�D�Q�V�����m�*�g�@��b�����7���aȻ��;�?�8�n��$v���k7�����o�î����W�=��4
9�T�,��y�i�@��f}N]�?�\�h�d���k��16����0E
	�e6_����\)p��Cc�x�3 ��j����D�DE�Dn���<�;�bd�ڻ�h34�8]{�+���Q��x�W�I�13	#.շ�����b����j��-K�uU�w�Oڹ�U
^~�å����K>�Qd���-� ��[��_^��}W>�$E��ap�G�R�d���T.���H�,��t8H���R"��|+��)�ϐ�5�;c�Y0��56�\>���"���#�������6���o�XP�ΖdXA�  �fU���N!=�����=������΍��!ꇹ�rghp��uuYm\T�>�;������:vշ��v�h��G��!C�r�.����R: )�����Egi�Wn[�)SR:!S��jp@�լ���;���>9|�&9�t���v��ҝ�[�rXB��"`#�������"�x��7�:!��k�¬�R�������9����H�h��QF����3��M�t:7�bv%r�.7мܾR긾3�ߤ�]��1|�FK#��%,�?#j���{?d�QM��e=~��@Seƪ&�1��dl����V���y㡖A?�ğ]����
��C�������0�a���[����}ƓO����?��n����K�u��+�J&����F��������Xlt={�S �.�e�ٲ���z�F(�xϒ��		H-Z|��sy`�����ܽa#����8�A�bTS,pd6�x_�$��l�Ɓ=
;�o���ԟ1?�V �~�U	��j�v2�a�)��-}�'nU��r��USK�y�C��N�� ���>rGώ�m���Nx�$���KD��4{R�"<���Od��`d8VI|��W��M���v:�Y���n�.`?O7v0��p�n߽<��P�43��F��+�W> 4�,�*G�ӣd��6\�{��;:�1��d��쿦�z�#@b�6����J� ���K-{�����M:�A:<w�r"㌛~O^~�}�!�䜏Ҹ�\����`�bDt��o�����)(%��(<9�a%�;W���02�7�ǜW
p��^MDk��|J����e��ݼ<�H�D�q�Aaa���߂��{k�C=\آ*����Dе`�DH �J����q(2o̴�9�0"P�S����{��n���Z�z��3,��Rkl�/�����2),�M��ֵ7��2_� �G`[���J�Qa�����(@)��JB��Uy��������W�z�����åu��q��Po��睍��rvN��}}��ã��C& ���-Af�H��tr���O��v����=�}>թ����;]R��t|ZY�"Ȅ\�d������?;Yb�c�Il��>���0���>ƨ[^���r��25>��]���?XM��-�S��~����sXf������&f�+���_�<��40}:N���}����Bå	/����}����K��A���oh��wn�5�Ya�3ɑ���më+1]���>�X>�"�0�лc�d�,�	SSP�y�������Y�L����X홓|v0��|i(�� �>b�g�W�ȋ��^�m3%R��I�B#�FIB��PR�YH&*sڝ�'n�	ݑ�9>�*s<̂F@�Lq�y�$��~p�uR�]f�`�6����_!����d	���}�{==�6n����}��r_D��n��NmHꮇ�z�fCn	��y���-L��T&�Wbb񚬽��
k��fq[6��46���#��!���T�������@"�`�� �� ,��6�\���	aL\�������B���5������~e7$K�K\"�Z��n\�̗Eڊ]\?k�[�I�2�y)J�4e�X7����=�����Y9��\�3E�͂��W�|��{�n��j\	Q����)LW����D-�L�E!��!T�F� g7��]��O��c�a����]g8<�JB�b����O�����Nṇ`L+��˗�HƢZ��a\����\BAr,�����"Dy�ZÇ?,����3n
&�g<�k£��A�{✹EƠ���s�74v��D*��ړM�lᅫȡ'������Sp ??�|�w�̀I�T1ds�r�a����� Z~��*�<�p� ��sx=�.
9�}~ Om$��"��"�$wv!s�h�A�r�W�7���|E��Îl>ey%n�2�2�9$��H3����ˆE�_�>��?N�i��N̈́�
�z'�>�H�䀘!*y~X��T� g�i�W�$���{}�@n1�T�XY�R��&�ۏ&���n�hD�� 1�e���c�
���M�ġ{��\L"!��� �����ņc��h�AY�d&A��[����ކ%�S��c%�蒰����NU�{h ���y�����7Ѡ��x�"P��=��8��?V�RA5��(���N�P���)�B
��v��w��U�7� a:�`�ì��ހ��~\���:ðax�V��!B�c��w�I�����FU��?[��*r./tL���42@^�7���8�����~Z^VA���3�A�Ie{
8�V25�*/oZ1p��}��;��6[�����	Y�����Y� ����Gb��L�#I�t'e/9��/��ގ�q;�胼d!�bN�K�2�̚F���c�F���f�v�w�ө�[�D{/M��4��Y�����X: '�����R82�_����u������ϊ�5OV�
x���r��ת���z̬ɭ�0bm�Y%��W�\���g���B	67�y�Z�r�8���2�O�����N,!�7�ukh�>�d�f��5V�8DM$���aÝ���haa���C�M�hav���w��ֺu�R#���i�Y4�=Ɏ�/���?��XFnor�x��r���l<�Ή��|�M����MɋB�<�?>���8��D̳�k;� ��vR�!���p=�+0F����`��X$����L���ӈJ��ۙ�0m�Xj�>o�?<�A� �EuP�v,�d����ԙurqK��I6RcpE��ܐ��]�Hz�Q�+f�]��q�>�<����#w��w��L�s45v���&�IMO�hmV���gG^��������wx1�Վb�E���0��D�,��Ww���-�5��/7&����-?LR�XF��(�i7sV{ArP��b?�,ݬ},72�y<P�Ӆ�6G5Y1��=[Q�	��+x)h�B��MuҰ͌��{�<��W�q(���	uRc��IU�� q�%���^�#?��龀�~jVIʊ�� l`��Š�1�F��ꊞ���AV8��ږ G�E��I��1����B�&����҈/��ǅ?!�w��lE�����ɓ8 ����'p{����d�yh��Ï{B�l̓�{Uv�CY�*��8�3>.y���[WuQ��#�Ղ��/^��4���J�!���Z+��A�����I���a/ߙ�����R�l�e���>Q�����6��,F���m�h$��6�,ݘ��ш}v�j>�."��$p?�.D����%���;��m���=��T�䁻V�܅���V����:�JƢ)�G�U����e�=~E�����a�#���U�'��>q�NF�na,@��1�D�?6����z¸N �Tc%�U���g�poB�����ϱYA��V֓����ay)b�+�����W}�>j�U�/ʿK��4�!jGG�1��?;܄�ɑg��>!���� /j�'�&�p�ч{�z_����՞Y�M|E�|�ɺ	����K���N���Jq��g�$��p-��{�����(#1��S"�"-��Ü�^����,O�&#�N���z����j�!-����`��e�����W��=*�������%��|�1����k�W�����Xv���ʪd~ނ�-���A��$G櫉�y��]�����W���0*1t7����S{|���'YI��&C���|�H��y�y9���=�OΊ�tG=�aQ1�r�޷	b���a �e�'�c\�����u	'��I�%�ѱ!��
ǡ�ŒT�쇈����ʇ�Y�x6B̧����C�� !����+nPq>�V��U��V�N��m�~]Y����l��¿-�����փq�H鬩�V*��wcsӮQ>��/���\�&.�KXᔬ�h��28��z9�G��L���(;��p�{6�}f���J�P�D�_��q��n��T��~��j��w���PFy=�N�e:�R/)_�ald/i�t��[RQ�{�3gS˓_{:0��f��wP
KΠ�櫙��������<�f�|�7�ntDD������|�"��Z��%a������#<�s�
�EG!�
�#����k����LP��α\�]�B����vr��t���U#�c�h%K��U�.�Wg� �Ҥnw��C`I�b�qَ�����'�w5w�C��	���։��C�a'e�dL�&P�#��/�Z�CӣU��5R�db'��;S�P0\W�a6�^�*l�$�Yl}�$8Y2Z%�t��PeFI)9�$�z��$��}��a7.�}�`'E���M̿��|E���>��.�h��C�������N�����D'��ܧ���鏾�_�9�j�g�h���}�6��;�n��Ƈ��"�u.��w|!Z3��{ ��@�N��9?~"X$D���Z��Z�߆�*��T�a���� ��#Q�>�8s�UH�l\����>�H�ɒ�%�d��ߥ� ������?{�����<7D�jW��רCv#:���طi���)2���_R�oP���=����mnC��Q5��[�p����w��slWvE���3�]mο^]�� $�!n�mg��c���e/��j�\�|��yD,�+v}a7�^�=̄�������� 2�+��y�ÂM@Bss��f���:�����D�]�L��?O���mMur�e1�N� ��q���\k���f�#�j�E��E���TR�Pi&��\a��!���]B�.z'� ���9q�B/{]q.�=N& ��å=�����������_7���r�A��"�I���5���V��a�ǻ�lǴʘ�S���^�*�ȅ3����CP��}�8�/a��07�{��_i���&b��D4>�˜Z ֡�+���k�!������ř����QN��A�@T��	��"(�|�g�ͩ���;/щ�dԯ-�o䖒��H	���]�,��l
G����R(����Nd�������lI��,�P���x b#��'AE�09d�w���>M�y��,z�2��pl�>����EM���V@ęrqъ�ʶ�p��!&�P/�X��$$Y~��y>�W+���=E�+��o�N�grw�/��m�`g������Or�o~=����I;�9��7�)m��7�*�@��ߞ2W&q��"�h�o+�ׂ*j��c;���}�9M��7�x�5���<��N{㵰3כiOr�{9�]��e*�W�|N���9��_:�uq�����.щ���BQ�g�\���̠M`j��_�a`/���V�)������������GI�Q���������6\_o��!��eۖAY���x�����w����TMPx~���)�z�p����Q���FU�o��+�W������5,�9�<x��Lu����WQ��
��(�=B�:�����CN���������C�8��M>LA���rNv�3����bL��$W�oqe��7�-�]p1gf#�u����'7�L>s��ô�S�OͿO�[Ԥ��E�̑'�m�P��A���j2�_�[�"">��J �z.��8������h'��'̯{��.\��[sfi������4EW�%���N�ׄ��j�����M��P�㿮���"*�d���
�i8rU�`@� &5l:A��w�H0wB�뾨q䥾C��4�}� ̣I���Nl��-duY��d���5�g��oX�qf��SP����mY�$�4���#b������Ag�Ҡ����l@w��$���`&��v�LKSor�h�0��5���|��y��'nd�4��Ύs?h:��\��
w��ސ5>�?�N3���&9,�$�w]�W�5Z�
�JQzl����!��D�����������r��@��K@@$�9G@��Ff�+C��(3��`7�wnF�M9��6Hp(����R.�<5c� =o�"����$��gr���F��vȭ�x<J������2"���9��j[Y����3aC��ܮ&�&�(+�@��}����Ǎ��s��]��j��q@��oo?}NYm���� o��5r[}�oO8�݄����s�p��u�u�g	�$hK?��:������g��H^p�s1������R�*�Ն�M��!\�k�Jt�JD���$�*��pX�b�"�T����pt�uc:�A���w[-��trA����L�Uu�T�������l��N����Q�3���"{l���̍�k#��E.8����$㇙�eX�j{���K@��8^��1�x=Æ�%p�b�s�e��X�ݏ��%�����b�Fd�g�G$q%I��+-ڼ�gh��ѝB����=��ۦ�v�����-�zG��$��`���-�j�.��"����.���&wzWG�J�W�NJe`v���'���
���B8^nA�_�>K,E���R�jedk���)"Ög�Z4���qr@N�B1y� H�����R)>�"p���i$�8�j���H��Pg��@���{jw:*_�y��?�����뛚~Lv�C3��ݿ|�$��l�����1!����Ow�O@���t�!B���sw���IKaS��*�I���L@�"�k����ۃ1s�u8|���O{Ro�~��Js��q�ϔ�],4ū1H�:�#�E�
H���%/��I[�����g�9�֋�?@�r���?͓���SN���!L��E��z�p�3��oj�J�d�D(j�j8m+t��Hv 
��WU�ŵ� #��(��|�Ue7m��@���]Y���)j���p�o����LPYs��7�_m)?��$(�b�?$�v���n���j�H��l�˱+r�X+S]9�*�z�`#����6��i�U|��C-�a����?��c�L�^��T4K�_��]�9�%���>(����������;w�N0�1@��}��孧��L�i:fd��A\Q.�-J>L' �po��נ�)��(X��ߥ"���:m�������Yy�Ye>K'xՓZK���KY���#��]q�VN��E� ��;|�Rm�ޛ�:IYٳ݉���̊o�P@`�d'k��廛����rP���*$��>|蚜O�c#��E�C<0^�_*i^�c��:[j�]��\bD'�"%Xp? .*�H���8*U��+��Rfb�MG�å0���Ax4[M �G�A����2�h��P�~��HO���.\E��{��d��	[�&����#%�<�A�J�z8wmf��X!K�m�K[�%�/P'�qq��$��mw�a�[��)^��hm� ߭�<Ӷ��]�D�2��Ǚ̆��k�=���>Q��c��zX2�t� �j{��xnW�E�^���#�i�Ù���g<*9�X�xzO�B���b:�Bk%��V�WM���/�S��Hak}C� ꯗ|��YT�
�X�&\�G�ǪU�'7*�m887��P�-��a�کl��1vDr*=�t���#,��;��IՍ�8�{p��}8{��K3T>�o�����v�9�F1�/�I�Rx�A�v%�A>O��7C ;�?2���)3r선��(�oᄸ���NhN���?������������~1�l���S�h�/(!�4�0Զ����%I����e���v���j��dr���.
��5�DlG�x��&d�]���	��jY��ː��\R���3@�*Y�m��nU�  ���//����;'�<1;jT�
}P�������T8ٸc|��(�P^5����&߯m���z��C�(�2�e�R�c_�՟�n�,8E����@]a���g��B��ۻ��&�7R�|<��(��,�U�����ͮf�G �o�UYp�^V�cC��u�'+�^LƏ��#�c.�)��Ĩ4��ϞE�E����w����������wl���c�m�y�~���yz��^7�0*��8�������1�&��#��,Q�̊?����G�B�߷��{�k������M��M	�'hd�V�4�^p�nY@@&��������Tb�R4Qzob����+�Ih4��M�����CV�	QP����Z��E��^����ȈX��a��������3�
ب�a���|+1�O+=}5Y�e�L��"м��=��w�H��j�����^��{֙R�'g�%�'���u�m�N�c$	T�k�O��¥���p[ᓡ+�N�_�==��c|h��o����^f���+(]��U���w�l1���`pL�������3T��75�2#� � +q����b7�5ڷ[�����oG~��A d�5��ǿ(6�����{����ޜ�$Ώ�؀=�p�3�Yc
t�w5?e�h�
�ܼ�~�6u��KQxo�4nwНh $q����Pڻ7Z���`r���-��t�S_[N�*�<q��s>Q�����J���t�[@����svi3P�#+���6s�7���7%��b^_7'�8D1D��Lp=���Z���l�+9b*���Ԍ�L�h�츭n�H��k�U�<�<.��C21�x䆡�G������(��^�3�Y�$5�Vؿ5n�sL�?=~�!�~6�eFJA��l��ȳ%b:����?�rM��d�S���l��؍��@P��m0!��L�C���]��%.Lbb���΀#CE�M�{�b��¥�y��w�.$��0�R�EJ�ώ��WH�i;��`u�k�y�BW�d�Cb����JZ����nR�~D&�Ǽ%2"�����/�"�j���X�*m=�A��q%��V����@`�(u�o�������7�O	$��^����������߲	��(��6uo�o
6��k����խU/�4��,������$mU���\�F�2�����Cl�pB�D�V��Z�⸉��	�|!(��7 ����S#�"8q�FNBH���+&D'�)�3���{G#hE���������@��6{�i������5S��7
| X�p�R��
fȐ�=g C
��[��o��_���`"�{�.1)8���TH�DRӆ�Fڱ#V�m Q�_�	����s_=�us��� #�zI�A(���;��G���jSvz��M�������ט�2�$s �P}�|$�Q?o~	A/�Ql3ⶍnь6�������+9�^$o	�Ⱥ���Ժ\�p��<�<��[0��)?^�X6�6� ��eO��KKtӿ��'1|����F����T��FX	'�!��b�;��`&���)p��χH��o���������3��j�a8��=w�n�ͥ���s���t�O[̢���U�INS�Ї2�q�����.+B�����le������w��_�~l��h�\]=wS���m�������ÖOt���S{|��,����!��>�Q���y�H�Qֈҷ8Ǽ��O9��������E3�.�̿�h�ِ����`��*gw��k1��`�9��̡(���<�I���X��E�aOiv�r���G�[7��]%x��8ڎ�ɼ/�yE����M*��\778z�ȗ&c�1_�/��������a+��ji`6�LJ&7弪Of��'�r-=�����ǂ�RλR��~�5�B��rŃ]���؊�0򗬲��qk�Q�6��� h�V\޴��W7z�S��S��.wL��s��L`-��Jp��_�f����>�Pf)��Y?s��}](f �a�\���i�}{���]?U.�Ud���%������/����s쎌��p��}�4�$߶�|ܽ����`�b��1
��q�ڎ�P��� #�ţu�>\b���a�A� �F��f�*m��e��^+���\����KK��'3�"�z������L `z�i��G�q%
��2����"V��T=i>�8f�}�<|L��6�\�9Bl$�n?]4d1���DIt�*:D���4����`?�ۘ���j�GD1mq�U)Tu�G{݊ӯd�"�,���؋
}W�����!�?!vsJ/��Sҥ��]�|�"��.��>X�����6A}A�a$R�KG����j��"���T,�8?#��mV�,�"�Ӎ�F(8�򶌬(�C�ۭ��d��AO��[�K�P�wNg|������"���O/���E���#�6��z�>�H��-O������y�@�}���M�	^�����.��Js�NT�<N( �
~�?��m�~��z-��g���Ñ�O�T]@�O���9*�����@�A�S�%��NzM�vx��FM������~	��%xք-ȞcЂc��c���}܁irp��/�=EJ�$�x��kCSh��N�u����F`� �p4\t��9�K 0�bkw1�3�ٱ�j�A���]�6 �6�K��߮p���>�� ��5�/�A}5C���ߐ"ơ������|�r�Ò���%�=Ħ=ƛ.�2�[�����������ℭW�l��[��m�Վ��}/{���^�������pԂ�/��vV-��?�  �5��+��n��L�s�x�>�A$��0��fM󪮎��v2���)I7�G?�ѹ�-BO$�Q{��p���j�-Q�d>dy��n[9�����E*���W��N��j<��j�~��Ͻ	��@%������Vu���H=����њ�$�Ze�Y`q���k��"m�N4o��K��T�C�����$��{���q#��� V=�b����FI�+L����+&�5�S�>X8>/���5�3�ӿ�ϯc�N�t����c�ׁ,�/X��X�x�k�ݢ��]�%К��e���@B 
�ys��"�e)ẍq�'HD�J��\Ѷ2�~^0Ȩ�V�$v�
Z���+�ea�يK���$�tH�(���+AI������[�`�6�^�,�,����C��ZU��*R��u�-��ͭ��?I�&���7qJ�����]��?U�_ E$�s����o~C�\��z�z]/�Nk'�L(�y*���4*�y-����ͯ����H�����ї@"�ZW~d�#�ê�.���"	)�S����<=2V)�+��ʌ���N@�:���w\��dn��#��c!R6��G��~��R@�No5-�}���C$: H�:�����V�5�b�����23���;]�~/i�Z���1�����*BⰞ�� �d���lg��Ĳ�'�Y��ų�o ���>FFA#Sy��ٙ�������q�o[I�mX�DOq\�ҺJ�<�6�0�p:��B�S!h*]A��A,��fɇ��1r�i�������jIT�uO,���*�=�p_�&(�#�mg�dX�.Ca��M�O����gv���5�<qO�=�g��V��Ir-�i�m�ê>�-��`��aM���ˮ�&���w���0N���Zҡ��s����2{���N���q<�Ob�׬|���ҫ�橳HvRs?GX
8x=�A�CK��c�G-Y��C�O<�H�*P!_�!�&���n^���Я:��HB ������ �H֚���W#�˻���:�����$K5�A��$Xh��ڠ���c_4"P�c�\,Kvۤ��醗�n��^�ﳚ��\{��	�K�7/�����;��'-u��u;���@W2e��!�����w�f�������Z0Y+a�u>��ZN���o��J[��7[�H��_��]��4��y�9�=�6����{�Ny�
����dY/	�� i/W����ä����q�R�Z
>a���[�<��J)��RTkݯ���e �ø�r�v�O.ms��/p�L�yO��h�|SZ:�!�0d�f�}޻��L����f�To���ݲ�x/o��|�
���<��˭�̙�jq��L�=B>!(	��gwn��`p�p2�k��}�I��n�{�I��4���sS�`�����������a<Nf�L~y銩
yoy����0�"o��&#_�`{����	��&H,�L���j�������S"K�=�cx{1�@�r�e����JX'��q���^7��T���k|�J��t����6zo�s��Um>~:���3�'f$�@��H�e�ڥ�:�L��Q��/��i�����OO�r١�ʑ��|�����˂�$�j���z���k�x�s�/ݮ����Q�����ؚ�F�[�R(-%��A�u���{�X���P*��ƖWw��Pďa	�@W��R����^9W� "r�`Y.�>�x����߳7��-��4T��e�p4V�����c.@bq怳R�X���F/-[���)�- �."T)�>t~���j6�q�]=����S�:�M/���Λ����`�2���&T�gw1���u5r��
r�f�ز�jx���xx\RdO^]��|0�1�;�-��'8��o�#�E�����h�.L���* �F���ѱ4�c�B�b��w�	��ߩ ����G�QL��.��h��u���T���L���0�N[l�՘6�R�+�>�x���A@�D�.&dw���T�rN4����@�tߠ��eN�F��~���R�"�Pq	h�}v��g_����d�~�e�\� ��.B�5$F�|'F���ϫ�!ɒJQ�1M(h-����f��^2����.Y��NO��տ-�M�U�(�
`G���r�B���o�f�T ���j��gT+*��"�MM� ����k������q;�Z������H����t�PK�,���J��+�co�P3��5����M���^�\��.p*�m27�0���&��ً�GG����a">^�2R�W�Z�>v�6j��������_�l:鸉�n��@ 'O�7�R��!j���8_�l���t�4،|�#�`����5���5�0�x��}�/�N0�O���_Ȱ�^�Kqx6�t"G��q.;��JB]r�<L���w����6�g���`B����M(�
;"cy,���Ǐ#'�������iI8�z�x!N(��O�v����#�`�p��֗�o��^���ؠP�~�ς�Z�F����;�4O�2Ty�v��K�����-���Q,�Ͼ\#����;�ty���7"�|F�x	���^��74Z���^��&Mx�H}�WA5�P	f�L�=p��B�9C������ꪸ��
w`Г�Hc����U!�$�Qz�#Í	�Rg��~^E�o�Pt��K:r��-��^7�b�y!g��A*sG���R_j�E��Eѻ"
��r��0�8L:]�X�L
���3��D���R`�p��ף���W]��>;MHG"e�p4}��0���z�i�V�`�iڑ�Gd�6.�ދ��B-���"�J>h�����<���e��b� )��~�1uɥͭ]���s��
,e�h_��Vj� ����	��d5������}�<��NT��es��Z��k�58����.G"<��%���?��]����x��~�72�"��o���`{�7���� �
j�������-�A)��Srz��}>�����p?SVټ��6ç�����-�o�[�>ő,�q.��à�/Tس�X�3R��!Ζ�@i����Ŗ<ߎ���X�u��sdl�u^�p'0�X����cL�Xt��mO"�`�]&�x������MJ�d���ep>��TֿG��,��g���]��@-r
�e:���Q�`�L����H��.A�������1O٤�M�n�
8��Y�,9x��� s
���
�,���8�h : 15�8�Ts��,bn���ǟ��H�b���p� �3���ĸ�����q��K��`�U}����j��Zf�̎=�Rh�j;`Ä�P[�o�1-J���9V�����������t�����H�M����<�6N"�\��_0a���:cSo���� �3�r4|��\�(��q(�Q?$�b�6�;�,Lv�da5S&ڝ��v�)6S
�8�M�z ����5b8��nm$�ʾ_�6�J��aE$� �L&X�vB(��c �8ٔ����$�=������k���Ԓ弻:6�i�*�Y�jE���i1Rd�f]!Qd
��-D�l��`���ρ�:>�
wI��˄��{Y7S��S��-(=�;�_y�Fp����2,�e������]�ww��@����Cpw���Π�9��{����յj�Tu���|ָ���Prצ^��Z:p��c� ��C��ߘ��z�,����C�A���>��I������n�y�Z�LKEFKI�-�.����Mџ��(�H�����ǫ7�GJ�{� *�����wq�����+���=�'���ԓdH0�
��Mӻ���m�t	���R�k����
���I�E�xr)��2���C '��R��|�	��u���P}!�E�#e����FQ�),jB_i�7���-����R[�lS�\�(��D����~�;�>dk~9���s~�a7a��[��3���l�bŗHSd
�ִ���F�SD.*<:@�|x����b��`Z�I%r�� �SY}����.�U}L��y��V����j,��^�
���J���	pc��^#�M���7c��`�ɺ��OL���8Z/�ѷ���.��ݱ���Cn�B�m��l��J.Ҹ��B��'���� _c��O?��	>��Q�-�+�����(6,��*EH��߰���w_-;eo��O���??�л�i?���XA|���#͝��bEL"<�XH�i������Y�0ҡ{�ɦ^)Y����f�>��5 �=��XinN#�!�,���.�
��)�N�_��v3�!�"�$T�v����@�-j|5B6�IEA}�����ف�������j��'Lh(C����$����FY�⥆�߷+X$��ӗ&�"��[�r敻�3��B�~�4��/���C8:W.G݆ސ�r_��xg���|GY>�i�8r�)#��A����=d�[U���39~��Ԯ�w��W���0[���.����H��*�u+�-�zZ�z~�
G�[�I�Q��8��5h���ӻR
ʲ��{��rg�bL�5O�������+)���Z+i}�s�5w+�p��_�C�}���2
�n��DɕQ��L�.y �_�����+yv�^��jl�~-E��& ]�q��=�\7(;�j���Lec��!�EL���-ȍH� ����H�&�ϊF��_vs{--0IS�?�w����:�+?�k5�&�8�|�O�o�Xh{v�`5��p*0�uf6��f9_�;�\Z�3����:�������9��t���\�t�zn�R�\L��h��l/3Ϭ|�&�� =���9��l�]�`�(�P�w�F�KG��dL�Ҽ�Yz2rK�����)������ �Wz�cC���/21�y�����T��<��kG�6�ʈ����������!�d�3ٌ��X)�B�Qf�>Cm��1C)��}�h=(Zm����- ���&Bu�Ǌ�)�ϛ���x�xW->��3��T/��z�}?Jdh�cEԮ���@ߚ	�Uw�iӺn�\}!�db�����xRR�jJ�I8MA # `�m/���7*���V�Z�F��&I[ӕ��;郗
�E���8����P�
ь�!X�u6��Z���C)(�	|�o�漌C�	^JQ�C�>- �񀏄�8f,[��}�E!B�Bd�FD�*�b��} �H߃"~�-B��\��7�o�R\.�-bξ��󃍛������;���\}p��w;o;��A�0�2�U�UM�D�����i�҄�>f����������r��n!��߰R��=��t6�������8y1�@����h7[qJ6��z$�<���DBGم�.�>O�˲kw���+UWkyk[�鲎␃1jEДΟ��%�"����q��0�2	*A�5ܹjP�0�F�Vi�b���󎵾�[-uw�^�8:�_y������0(����,��	[�Ȝ����)�ehe�i4�z%��x(w�xym�Y����t"�Zq'�~�^���g�� ��B���,v��D�W�h�,�ǈ�U���W�7���$f���Kۑ3�k��J����x�x�������^b0U�c�	ɇ�ⷷӨ�d�E�=�l�L��w�, ���G�0$�4zn���{�4�)��.}4��z�ۗ��kw�p��j�)������l� ��*���յ��:L����Q���пRbҠ/:��\+PE>��d�VԂ;Y��ꁋ�����ϙ/�i��brk��
�]�C}�y�5U�Vc�k�Yxh(��Lv�*��߯�s��V ]�� �� K�m��#t���Fg��b�=���\e�S�n�'�誉�v�4t�n��&N�IO�����B�ЁoJk�U�5><�h�É~�+����njK�lQ���ξr���7p
��OPO���Nٞ7i��<�����8O���&D��tS�v���\-"��48<ˁ"�&H��L7�1��ߤ�|�����RlP������*�A�C��F|��}����#X�h0 �j��|wcI�sF����UG�Mg'���x��j�a�חh8C�/@Az�Qcv����JZb��t��Ϩ�+�{܀Q�X�C� =慤Eb��{v�g_e�jĔg{S�T���^�%��>JCV�Z�(�{�Q�Q��?��9�S�t>��T����1a��m�v���Sms���4�����9}K��9�Ё�X��fw�ZX[�y q_�-TЭ�h����ğ{��ױ�^�b���a��u�t� ��!�.�}��j��t�]�3�"�~9*�@�o1�X��S:�k��t���s�@��e�H��8�/���a��Dk�2���['/�^ӊQ���b�AV.�:3ı��;
�=���Q�*�9�����UV�^ج}�0�#����q�k��:�?n�_y�{���-�δ[iC����	�Z.(wd��m�H���E ������k��C��ӫ�'�[2E���U=.�M.s�Z"�{�@"�)��΃���7�8wbP��#�M{_� �)�o�v��x��؜��E�	݋�SFo�x���<h'���:����)M�9�J�2��4���b�2I�mQ�F�Z욨��"w脸d��۲���<���y z���R	�����gu���-���0��g�;���FBfj�ո��������3�X��R"d�m=e7�t4RE�[���?2铵���?��E�T���_C�U�#�|V�~��'G�2b|��ҶAN$*J�(m���R���-�����	�'AG���+g�^�P�	���� j-����~�o�>�*Pr���o�e�"`d��yF�m�x7�z���u�HX�)c��Z~������aO|�$$3�
��O��͙��K,��V���>r� �@�1cc�����u�i�l�\�ڞ!�UY<�K ��&�roj�X]{9*�
Ð�n��3霕2������EQ�|@ 3W �;�2��>�\�����|�}<mD�0���1�'t��� Z��t-f	�ڏ=��v2s�ŲX$���_��22I�;�j!���b�	\�"�5�|��!����ʗm	�w8� ʍ`6W�4�?�n�棶���?e�+Z���;��)��A�t|�I"MD�#���M�-\���?_E��9p��@���<GB����}�͠��Tw��o�['vW*q�w䞧0Q�	6ẄIiL�vv���>w��%\� �P�R\��D�����q�B��R�[��}#��߉�~�����������M�k�L������~R5�B�-��
ϥ~/:TVM�i�8�r�;FaԀ���]����IFJT9�)�W�O�o�4X@�-1�Ly_d9�+��2L7YV�U�K�8Ӎ��������C�����SX:U$Ou^=�k��%hg0l���F���-{#W����@NOTLg~LT�>�$���J4��������ZȚ��'�V� ����!�<�f&c[o��7b�2K��ˉ|� ����jH
� <ޠ0�F#M��:�pV���ܐ`Ϯ�� A	%}e��u%�l���+����;M_R��D	���KjA��I�4����߫	�ž�2�K�#+�_��}�mE���H�̸X&b���ܗGi2�K���$��<Ī��3�i��Џ�JK�S�����U�%d����X0,���x3�"P#<	�15U`H��7{Y������zn����J����!y��b���(�~��b�Э�}�\*��t�������[iLM$�M^��I1��� ��6/�Q�1�ÃN����(�fo���k�Զ�)]"h��w��_�u��nR���3��Eti����f(��Dy�ŪZ ����k����l�q�+�s��������褦�U8��:9�x��H$w�xexc���GX�k�����̙��V�lX���E��%/Xp
mm���=���[�o�>H)�b�Lָ�8�Ų����p~?-�RF���?6���Y���)���nP,��B�ʇ���ngj^�</�]
ʺ�aa
�k�@�w��2/��7W�M�����L�:آ���p�ʆϛ$�}[	*Gi�t�+��YE9���O�>��!"�q��[����e�ڽǂ!��D��K`�������0���ހ��O��X�Q�F�L���$�Seb��9�p �CP�w���ꌜ������v7s�O��au�kꍻ<��6RN��%2o�nnd��"���%+s)X�S�u��F7�j%�$��W{�W��T��:�`�5p\~not����h� �Z�I=�:u�[�8W�<]�]�cS0L-�T�B�uP�mu�u/w�o�뀮M��s�P����[�F�x��~;jMG?����-��{��-'A8��j�Q�>)w����W#JW��\̀PN�O�Y��$�쌈�=,���Q��}R�FCk����/�@,Xus��s'�%7��D�?;6�C��%	4	�I�\��`S�H�*M�@Nb��x�U�_�9J�IDYy���uO��駽�[���G:��rE�����WW�gh&�C!Y��������V�{�M�"���$^Z�+���mM_P�)��:Rik_H[>����r�*�?��6Ń�R!dzq���{�"�q���S{{9�~lII�<����_x��t-�yO^Nb4[\��sc��B�.6�~����W����E��M��o�=ۦ�p�3n�Ǭoo�$B/��pi�Vy�ï5�d��*�O�}+�rx�@i�-�O�T٫�FJ줪����_L��
����p��N0����=��PR ��@"f�vü����9�>t�5�pvz�g��Z���b�l����^��E@5[I�_�MP��=�CW�?�D	_y�G���]�a�?W���O�A�}�N<��^K��@q}yƣC����L�*�b��$[R���y=;SPN��ay(���P�[M^:�=�\�)����@�w��B�<

c��]  n�"a��y��{b�_Պ�J��F�ͪԒoE���:zk�x�6{�=�{a��j�����%���<�^�O�)(q��.���O R��3<H� y���nM���m��]�~iŅh/9�+I-,�:�a���f��B�"�3���$��k�,���,��9���=��]�?:����DGKkm�j�!`%�B��H�p�V��IjۭjS�L�ށ6����(���~�����ڕ��h�n���B�e���oG9�d: 4�=_�����d�"�AaRm�=��%�M�0����Ҋ�6\�
�7���d�^�7��Ċ�Ȗ�� ~ � |�P��\�.�"n`Y���Y<�x2¶.����+�|�ɴ��}�e���ѱ���LMp��k2J� `:qZ"s��E�X��M.a-y����x�\�7=me�.���ǖ~Iwn���S��˿��*�*�=*�G�T5�|sS��'sNLr��}��ZC�bλA�S�
�G4 ����tg�� N-{ޞb��Dd�j^�
��rHl|�jӦ�/�M��>AF���lEm�-9:�Bg��`����Ţ<��H>��$<��։�#�p��m��&��Z��<�w5A���R=қw�iyn�2��5DC��E��
�E&������A�%����7 ���FB�[�|�j�����w�
�3�{EF/������j+�� ����`�AL�	kEEȵG���ʔ��ۨ�k�*-�h�j�Az3V��rr�4�r�)%lp.'�|�Q�?֌���e�6�brmI���]�<�%�A��7;�rݔY,��x��5�ٽe|���%ް�궍p�Br�n��0}�'}��(ϵ�"M��y���3�i��Zm{y<��ğ��/g��뺓��y���H�]�.�d�e��r�&�fL9�,zxQS���onL)�.R�q��>m�c״������1@��U����M��M��G�.�lp|�P�����ك�h�f��E�� �xY���������G�f�����E6ڒ��poz�3ͫd��`));��,z��!/X� :׾����}%��b)E�
���{7v~�n����9�}�#To����S��n�����2����o���+a�+�P�/z�'6��Rt�x��%�C&b�og�u�r�@�އ� �%'듞AN�f;5VE�5_#z�;�9��6����O�B������Ww���RE���l����EɈ�Bc+I�'������r?�}Ӎi����дǈ?%aj��M��>n�&��<f�Ǩ��G2ÊDj�	�D���:ɪ�ث�%y3����Z@�͛k���#Pt���x�=����<%I�诋llN>='6〦D1Ѿ�������^)�Cw��_�e�5�Z���V����{��S5��Ϡ��ʝ�2�����O�]'�������^2�������Ca��ᨸlf�*��X�A���=�����;�P�T��q����g������V��T�/eM���W!���BXϥ����x�4,9ۄŷ����dA$��id9x�q�	)`������]�jG>�'*�]�t�K)��KO'VuWvUەv�(=�����_����-R%N��X���"��ٗ44!G��3U��S�FS;ʧ2��աIឬS�9��o+��jf&z�i�lo(��X�$�7�@}���^�p�'���c�AxIgArJvHXϵ���Շ��u��0}�]s���%'el����a.���T_�<w�~��J��[�;j����-����7�"b�u�VZ���+*��-G����x�U���+�.�=����~���;���v��@�W^u0�(�@Ď�kL�LG��s��:��LIB
�tu��W�j�8UQF�;o���c̮�M��sd��<i�H�`2�6+����Ӥ]A��i�X㟹퓣_�I�����6�v�~k�^,�����T��8�9��cd娌�%�d��zDU,�x���O����#��Bc�	�q��~�.��,���_?}�RH�/�Ϥ K��:;��)c�]�p����@OY�5{�t����;�2�!�����߀n�W94��-�|����y��-�siHEm�,���'�*x����HKH�^Wjeq ��hV3f۳l���r���-,]ŕS*�"u_�D�!��üx �h��*���٩��Ҵq)���4�ЭY�"ȝ�� �W���D��[���`H{�0��&���(�'���O�iɭ"<��-�K���%�����=[W�!^bS����!�y�c(t\�D��Ǜ����o�e��dJ�ru���/�9A��C'�*��<���8�\ٛ�� I�.;}���?��N8�J��
.�]����J���-s�/`%��+:�^[B,�_h�+�ލ:?m�}!��0���Ig��~˟�����-�.�S~o��,`O�O�˾�-��h���h�S����V���&M���SsZ���)�A�|3<.�sb�R�S��׈q��ӂq���5%5�&KnqB�(${�A�6�K�]TQ>�������_=���4#�r��5u�@���r85Bg'�(`�C�D�v�ܖ�6+X������|���=JIns��Y���DV$�vr���	/��Z?F�h�da���G��c��eS���i�da昅/E��KnU��3�M��>���I�H�{W����
���(g�B�cp�df�0kd���a�����=e?�D�^uz��I7��{����h@��gٳR4��+�������2��S�9 ��tzK}��>�0T���Rz&�f;����o$�C1A���ֳ��H8�<w;��^<e����v��H��A����x/+m6K
:=�wq��DNԄo(
��e��&���-��L���Gp���2���u��1T1&�Xm�g����_��|�{i'ȓ�2.�D��x2a�l�?����}XZ��#��G����v�aZ��6�ؾ��J�)���9�{m��Z��i�����A�ø�]^~���)�Wz�cvj���s���垱h��r�H��O��~��� .�@D�(���z��v���ɠ�Hijx����։��w0cf[�~�Lw	���`a��J�(�M�e#�ɀ��S�G�b3H3@����3�zLI�~���/����
-kj�^p|mvd�gIO���\&��Ѵ����T�W�l��,b<G��g��F��0�0���<'�N��8P�{��sm{���ٱG`5ԭ1l��g�&%����U�^�-uLII�,���J�����4����o��͋"�G�l��5p�C1���>�����"Tu�Z?e�,7��1�0V�/T5�VR
�FEa��~�������-Ծ]+.ꓐP'f��N�Dw��������!,��-����ex�Q&)-?F��O�* ��P]?c{��j��l� <m7Gt#�L��G����c�؟�	$hH�H!ڗ����w��69�W�Ȣ0���_H&�ަ���"���b�H��L�+�'빻���gJ��8^�G^;t�j����{	J;��7���� Ot*n,� �֖үH�@޶�M�@@4�éX�.Xܾ�?�N��l+s���^��	d>8���6��?��HR�sB-j�Y�V�u�B����D��%��,��T��*����X�x������r�/b���^��S�Q���4�?PK   ��X�䓶� � /   images/132fbcdf-34e4-44dc-827d-09a965026955.png�wT�Y�/��QgPA�H�%PP�tA@zE�&]���E��@�H��~����ݵ~޻�]�����9g����}�9񉸡�u�����赫 G�#'/:�f`�(���5�C�:t�1����z���k �w������)?3?COG?�m�u�p����� ���JS:�@�E\��/�{i SB����[�?���s�?���s�?���s�?�����
c����A��?���s�?���s�?���s�?���s�?1..l������c����DQ�;1����9[%����-���w}��.'��3;�\�/|���Wh��ж�w���t�i�%��_��������~�j��w����P��S��OZB�v�3r�r��E�8:`7�h֤���`b�\�o��{"?���s�?���s���Fq�� t�t�k��iWg%��ZQ���X���9�G���N�Z����谥#�鏀7z7�;��]n[�PQ蚭0B⏣��/���t��/wetiD\B2�Z�QF�:�+auY��f\�@�;j����+������'F��~ӣ�+�qͪɱ����E$��@k�]�R���.#}��J׽��L:�Ʌ�?/ZE(W�A�*�>��,�gT��.���V��`/�Y6�l���g��G4��乄��6K�E�k5�	/��u��]TfTz�MDڝ�==����D��T��y���
��=���]��|�	e�i�f���k�N�O2"����2hە�,^�S�Y@�&���2zf��K���y�ۻm�ʵ ���sm���Ȅ�WT�J�=~�	Jqi���.��g���r�u�&����&�+
2"��u�����}�۫����<g��:��sB��?����
�m݁k֢�97�����F����KؑQZ��v��6?QTj�M��	thf*k��}H���C��ߦ������^0����hKR��AKC{�{|]9��3j{4��������Ur�t[Uǣsml��o߿l<���"Vi<H���xb�lr>%G'�+�`]�h�O��6�rq�3
�gbxN�\��il� 8�Kb�iՎez�����N�]{�Ҕ�-I��m-�dTy<,5PF�ɹ�hX�o���md�^���s{ç��~��~�,|��; a�i�7#��ċ�SB��:�.b�vUrs��Um�c�ٹn��I4/"�Y���l��0��&�U�ptY�MY9����T����v{�ڞ�}O|�H']�qA?�.#)~�J�.}�n���F�H��H����S�u�O�}�)u��Ӫ8a��{��%����;����m��k��SK���ɺ�sYw0�������,DsUz�l%�
��ʒ��q�G�1釠��``��m}��Zz����k)%i�򣰺��;�M�u�*�/W����z���I%1ԭ`�@��y��䪧�7�SmƮ�u����u[���\��G�Ud�ב�ڞxݎ�4l��M屵����{�w�h,�b���Zzc؝]��	�#����Q:)��	��^d��Gv7�����I!�q
��>������ƞ� ��`0�Z�-��%���F��ڒd=�,Rm��WvG�A
M?W����O��/�;����-U� �����x����ǲ�^ 7%b)޷R{:r]<��N_ ^�}a���� ����Xw��>Մ׌��2I΁/]X1"g�2���@΀�jU�ۄK�"�l��Urn4�&(�&���/V�����K�[�����7��>��D���B븹C&�/�٦(ԢO1jk����P7��Z���봵IN�����v�:I������mEZ5�=�3�b2�߃��g��p�����Hp?M:��9����v��;b��Qw�Rz�D�,c�J����wF5�z�sʪFW�}�ޢ2z���`�̬�J4Z�(�2�r<.�&��K \R���>u����is��U���O��J� ���Jޱ������!<o�KVI��\�9���/�1UF{Z���=-1"�)�H���h�P�F(�ȥ�L	lB�i�d�bՑЂ)��1����#��~r�����5s�/L*�$�}YI��l̵Q߀I�o�4�2>��IXjھ���x����p4��᲼���$$��7���i���s��\h�o���ڤDBC�ս�d�u��u"Q��4(�_#�U�4���˺��2O�s�A��V���ᗛ݇#d��+l3���pC��̮sc2TE68�Iq�BD_@e�Y��I����-�@�H/��
s��7�~1]��s%��d23�)ol�v�֏��)"f�l�o��3��������jD��Q~C�i#��#�Z�4���������F0�G�1cط��6����VeX�;��>��>fy��Z�v���|¹���7�d����#�
��d=�2��~ߵ�Ξ��L�U��5���O�����ۇ+���#v-�TM�/L�&�V��ѥ�޷tB���[�mh�9��V���D����\��|D��v�X'~�1�πY ���)����� ]q?�Ӕ�����<�6)�xz������Z��UlQHG�y�j���� �G �IH�/�
��5�@��b"M/y����7M���a}<g�VY=7_7�`���&�b>`��e�P~�Cy�lm.]}��K]�}6Pt�V��"#筬vr�;�\���T�UȜ�� ��C;H���T���r઴fQ�js��&�V��y�e�-�G�`d�H�l��8
N-ib�����pK���S�Sݳ<y��mo�u�� �LN����2m�d��4�WR�w�<�azcc+���gz���u������V�e����.9xy��u��A-�&?U�U��j{(r�D^Nx���f�7�$���u�LȠ.�~㘱���ҽ<�Cg���'B�^Zz�;�=���S���E�U�A�O��*�Jn��<��a�?�ܐ? 㿯�V0��kq=:Sr95���h��-nԘ>^6����:�J���4G�����%�u<���
Y'�=޳F�u:�z���%���U)[�/�{�*���V|��>�4�e3Rrx�K������j1| TDH��dx�+XfP*3M�,X (�`+�2$ X�f+��pE�zf �������Z 6�xx)������A|�[JUN]�.?ʯ�3�>쏣ו<�p�v?;�c�dI��U�Cbg�L�����1�Q��3;��]�+�_�],`�;ژ�Ņ)pu"�E{P���j���5~4��GѿC�A=:r�q�t7dwz���{�E�ȸ����<��_-�Лo��׏%�4��8mD���>��{%�ш$Id�[�eYk0�m猧d;�t;B*��>[y�-��rD��[�ab:˟�ܨ��|�x#pu7������}��m��=�5�Y�
���|f��5<�YL�L��TbA������u���E�I�U�A�9��w�SlM�3wI�����L��������S��qU�ɞ��ۛ�x�L0O��T����}j#)ֽ�`�:N�ҵ(��\5��Y��um�=�"�I��J�|ro.{�"4�
rI}�����ux�Ln���[�q��g���/�u��\I��ғVY�Q���K�!w�2�yre\X��'���B�*d����"����ȼ�*!F�AΨ�8�B��鹻z�G�M;萉_���!��OL�������}��3���)0�Γ+gA<5����%�X=b��C��`��лk��=���[c��{��އ�X����f\O����~�Q�����0aru�*�f� N$�\.[zh�p�5��˫�E�Q��
�t�Ū�p�o���s�q�~��5N]{�Ŋx���b�ߢ�y��<��dԣ�j�_�G�������a�R�}�$c���5gD����������#;{�;���a�R\�o蕱��9����)�BBҏ$+���D�1�!�ĝ�8��T�1��|�Y+x3
��65���o@<\��,�0U�a�kJȔ��?�u���XTG�N��{m��
0ZH����U�6�Y�պ���&����b�&��\����y�y5����e"N2gK� k��0�xPҩ�/��]k�WYn�]��@m�E�^]ꍪ�~�Y�frF鄩�p��0&�;��{��ڸ����W8���6�R���bb�:�P�#6U��ms$A(N�o�6(nU���[{��&�<{�pV�3��W��$A�:' �0G�L��Ě� ����<��U;�6����z�d1N�8������A�ʃr�;1��s��E$|rMu�7W�y��P=������O�X��q�Kυ�'-��#�{�x�$��c���=M�b��MP�Flv����������ݬ����`]���'�Ω�s�V+D�5T�v���^��f����j%m����f�� �A�|>Ӿ��L���d��L��v" ���r��,_�f�Z��?O|��j���]z�����<�������w�!������n#�05��lo���6Q�^ǿ\xsP��^�I�4��xc�UG�A3�O�dݹj%�/���`�������(����ҕE��v�}��*��s�m��`���wz�/'^�N�!�p65G�˝��Fj_��s�E��w��ǫ���Q`�*e�r�>L@��VE�A�θS.��&��P �]���LT�e�Y8��O�)�I������8[}��,�Q6�.���.t��.&e}//�l��"��]5�	ZSIE"F�����D̨r�N̎/2��I%�"4��+]���c�Sv|�(0�ۏ5�U�M�ߦ�x��q��4��C�,��uEQ�x�&�¿�$V�&ۖ(�0Q��)U^��Fa��4�Tgu+���sC��ͳČ$5�Y`dY�|���U.{���X0�1�1�>�2�/zi��xl�I�M��G��Mh �_�\VG�,�D3ކx���ƣ�0����ZI?�'��J������F��Ѷ������իn��A]�E�4��j go�\�H:93yBBT�7��Zn��Pha#1�>���L�j(�*x��ڌ'��+TEQҹ��Uв����{-��0���g�m�O@̖,T���mE,=5�C6�(b ĉ�E��
��L��T�R?��M��V�|3��I��M\�UПZ�iTF�1��1�1^�'h�CZGl{e�,�1��,���^�d8 �u�A�$����N�G�αCl�ɮ��Sv?����˙�g�A�NX4�]���o�!��쌢�wYA������&��V~�܍�Q��`JϏ�nG���=#�lf�ٴ¶c�`w�X��� ��x�ӥ�<A�KOC��x�@,��#�s�vO��!�c�(V���r>����}� \U�;��d������j˾x�^:nv�xN���i�Gb�n�p&=2�}�(.�!7�����[ ���W%��!��zr��D��!��lm��Z�rr<Q�?��B����#���o��+�[�nA�}!�7@��b�>~�/mR��쵫������s�y���_�`-8à>��q�V����q���2����g�r�n>|��f����Ĺ!�BB�cm�	3r��kiǞ�\$��e���/�.*�1`TغJ}u|�Qa@�y?�̛��Y���� 2�F��|O�"�C��BRa�׾6X�aF9�oV��B������Ч��	��4��<T���W.��Z"D��\y�������ƍ߇�i��#Jz;�!4���h�}��E9��I"��
G}x����<�E��g,�0���A��
��.�SE������
�A�l�}�6g��ةS�uk��>�ghi�=+������>��k��c��|�Y��1#n��8��&�N�<<Oj�CC+9�+K�WXᜱ���R���>A}�B�<k^�W�qW�4$���'P��B�a7�q·[�A2<�����VSѐ��z�B[�V2{sȢ���|�n!���p��)/&���ΑU�W���w�6��_u�E��]�\���O	����)�-���I�B�y�́_sԮF��)5_���9��ܢV��sͼ2��˖�U��U�>��dX?9S�����F *���'��:
lg!;눻����G�B�������W���쾿���H�sV�A�/�o�Q���MI�=����J!�tWl�U������F��&�y�A�NB:��%�Tf�#��5�-"�����^��_��z���@����!l�F�'�(�X�K�1*��ދ��dN=z�p}�$wE��G�n��+��- ��0	�=��2j�Z,*�-z`�	ic�hzf��R�����om��^�����Q��=��8F��$bxE5+H�#*i��1���7o,��޴��s�6��]�ƻ�Wn铲���U;� �e@��-�͌u���(���ֱK��v�LV,rQ�rGE�$[	��<�7�k����N�ċ�myxn�.r��/b�6
rm��h�{I��'����|���W��%��}N)X��o��P�z��X-�:�1}���{�����A�iH�	��km�{���t�M�^A�D��A
��QNb�DO��Q<2������~I�����g�7��P_�N���E��x>���@i1��~:J�BU>��K�\.�(�"��ē|e�^c���@�� dS������4�3�{�'�<k��=/�>$Z�AQ�-������GĨ����P(������=�$���9V�qp�,�y���o~�]�)=����	 �ziC���u�7����J�~�JUE\M�T��Dq*j�^ �~�N��T�5�L���O��1+K|[�x�s:�Dm�My;�W�����~;��	�zO�Ჺ����!�2�bc(Fq]�<b���v��*!#_�ַ�҈%��]P> �E3h�MT�
^8��ӳ�~�6g'�#\��\g#�7������v1��������\�<SG�_[ۏvx��J���d7���_� 4lご4��.$��l��Wn���OhŜ��[V���a��gM
t2���%S�ĬF�A� ��Bo�|�[�{GN��߾i�~��2�I��_�"Q�N��}���^&uf@�W����� d�"�i�,���z��ؙ9N톀,�`�mF������I����o��l�4Tx��W1�M���?Cn��W�7����;z���T�glŜtH�ߝ��'C�!��?TP��C���������"
)<۶�1���4����y�^�v�yw~�t�ze�f�5�{!�Aslgc-�Ge���@)�ϡ-��z��*��8R�����Q9��[�Q������L�K��W�%u��}18��v@ա�hg��}{{�GyF�Q�Ql���7pc>��Z?Z���������(�\�|��$���5������wh�G6pg1P��8�c�?'�u[=�J9{��L	��I�-���ݭ��?rk{��܃nھ�X����@P�p#���޳SB�&�ˤU8�ؒ�?`=���Z�$�8F�|�=�⋠���	-Y����у�^���}$�u�ۊyj��yx-�`�Q���Lp�Q\*��@��aЄ��t?���jp��DNj$�LqV3,9�R���O݆��;3q�(��5������n�x�b:�!$�a���26����(J總,�=
�0'�ϋ���!+�TRPPWJ/�>��T�L��m�~@���jnI�݅{�4&D��
��ܔ��4�������$À�"}��q(� TAG��4��K˪���p���A,�o�\j���|�D/?�3���y��@>`��L�9�K+��W��Դ虬87�ڑI3�a����$}��
E�,�
o۷xŊ}�@F�X$@E.\��rf���R*�1���x���>���\�L�����RSM�Q���yOX����C]DlvL�M�s;���cW�p(�ݞ>,Bw�^�?=��+��%d��}ˠW�Z��k��Qx�3� ��o$U\]���u��l'/�D����VP*q�`�k�Z�ݓ��V���i�D��C�N,GJ����)����4��Z�ɏ.\�2H�j��I�.�S��h��5��M����ʃ�A�)s���읔��_��q�uC��q�8w���.xm[)pm�bpm�I]�~=w0jZ�t��e���`���A��A��~T�>��j
$�mYМ4#p�?�#rg��'��Yh�;Hj�eWd��w���W
6�{Rs�[�`?�AMy�#:6�lyB��� q�ի��}_��6�=܉���j+)��� �L坏����j�)ۼ���3;��Y��I��7$o��������ZicD �l���ksv���VjP��l��&F���pd�&AM��m���-MG��*�̏��B��N�v��F�9�M�C�	�#�~2�����CsH��Q>3b�PڎSna*LY���;ڮۂ���H���"��O���#���/��K�Y���*��P�W>���k��m}iCkH0\r���	w�:��ua�3`��k�w1�`�~�M�U���ـ�}�!��;�`9����Pw^�X7�[�LU׶���v�cKѽ�a����!tf�NYL#Yv�	Du��#�y����̭�_mF�`���
����ka�ƥ�W��	��dj���T���ؤ\�[��\�W��]Q��תv���ci�wh�!�@Y�d�B��LU���5Ņq��Pw�Z�ж��^���a.�*%� �Z���rߑ�n�����_l�?��x�x������o��b��u4{Z���v�����αQ�T����WN��W�&���ɛ��I^۷Ѽ�Z������OT@]$��[��0��K5�@a���ۂ[ƀ�v�0K�F�Ԙ��Ǜ���˗�H��Ru��s��DH��/�DR���9�F��jS�A�&Md�f{U��f�M�B@;B���؄܌<5�/���:�+Bѳ�B͙�zaB(&Bf�F�#gԅO4��Ze�]{�n�eM9N�ʁ=U=�uKc@,#>�n�l�H:����f�Ǩq	4m��>�g���=��K�yG�^�~eM���1��Y�w����^��7x��V�&�����'#�8��=������rSQTQ�6hs�eʓ�\m�����gi�=֜~Ec_c+^!C�݄��?S1�""1����U��l"� ��/ w��6��Kk��1\.�����%� ��#�j�#72�C|'��l�����M�-w"������7�0�����h�#���>_cc�7+�����T<��0կp���l��^�6ȼ�:�r��|�m��x)����{U�;ӗÌ�Ƃ��vJ$��ڟFo"�¹�n��H�[��`��S�@;��$M���Y�V3�cY^�|�X2�w��wْ��;�p;F��jo}M,2x��FuǺ�w�@�=<��Su|j2��R�M_A����Y����$e�%�/9v�6\<9���8��@�m�tY��2̺� xmGvGi�L�J$W�[�����6���&���Q��Anv}�S�pb�8m{`rO��\:�N$�nT?����w�i	�n7�O1��"�;h;�΅~5�>jj�[įJ�(��J��e�/��}ȓ��=nAC����).�wd�V���,�\ś�������4D�p�vB��аo?̟k ~1M�&
65c��C\@��K�.�R�郹�,1�H�r`F��J�,�O�����G���U3wgiB�L�v�D��\"P/�6��%�f7Sm��+Ӝ)��|�g&��qKި"L�?��4���u��r�>T�lu�b�У��=���WoS���M_�F/��KH���җ�6$���(`��a%#$�Sc��[;t���9�~E\1q�b��'�0����@�e��|c#�i�+�]k}����j��s�h�W��&�@�v9|��J�֜��P�gZ���V1[�٬#'}�G���R��}��ؘ~5�mȚcJC�<����9������b�~~-*������2�5���K�*c�X�=Z�R��س���3�����^�Q��"J�o��sV�V�b�����dB�e��_��ձ��,P�ٝ�T����w�����kaJbm�ѱA]i���hK��ظI~y��G��&0$�!ɤ�X���9��d|@�Mu�3��0��%�@�Ѐ���X��a�	�&����N�we��M8k��~�<
�PYj;������?��t�ϱ(!�}�H�4 l��{�x���Y`�j�;�=��C�<��wd���&�{�n���POM%6�#��q�>�0#1#4���:��!�X�0U|+�Lo���A��3���Σ"��3=�t�z� _ꔭ�\�;���L��k�3{��d%��,����@p�U��}k����w� ��o.!��8��ɦw`Zh��wؗ���W:���}�^����z�?���@��MŁ�I^2���P<^�IcB9��������w�"_�S!'S�8�7�����P��
�EO��\��xbuݰ+��qߚ��;�<聲[�w�VS���{��� �N�f�@Ƨ��Eu��qb��T-ǴD�݁�$1����T3c��!�V_�:t���4�c؟�9`��ÖlObN=/�5g�>�U�6�Č�Ȼ[R�^f�� �.���0�{�=�(A��Q��k}{XkN1��X��`��NU��h��0Y�f���]=��y��5GoM������x�
.�t��F�v��.�F���� �e)z@��\�&��ʼ�}'7-qv�)������*�u(;չ*7gh�AM.E�!-��Q}Zި���e޳;�Y,�۴ẽ�֋����|�}{N"J�7��-u��T��iO����q�u�96c��{�|��
�N�AHk��m�^�T�X�'���x�����0�"�M�a=���Wvk����'�q�k����Q�:�C��.���nh��zu~��z�z��h: �-[C��6��N�ǻ��a�`�l�_Ā�q�:���2�i�F�Y�K:�Z��S�4�6�_E����&W�k]��z��I���g��׭��[�`�=T
l;�g���֓5���ꤍ��r����n���4vٛʦ&��*4c���q[:K��/�G滑8�7�M��=���'�m7�K�A&o�Lu�I�S�o�4���&���(�J�r6���W��o�?v��@��iWY���$�Wty^���eo�/U ���@����Q�ٞpG�{�/&&���=[4G��\p*�p��1l�A�A_��2y�3�/շ����r�޳���������l��.�\�V@/��	����?�/���_�R�#�����'s��]�x��[? M�[U,�'�3�u3��&c�ga׹�j� ?�+y;G��_oR xg+����՞	���Cg.*�󒇛�,�i�1Vr!P��Js�>��^]ҫ�؟�ZC�[:�z]>�R�,�<t?�K�`��Q�^r�]��]N�N\���&%v8&���I:5��aw��Ƽ����fڑ��N�q����=��zN�|C��g��c��?ί���@��s8��~_x�n����kJFy��Z�3^��6@��S��U@��_l�%���.�l�m�-�=�l�	8#9g�lX�۱9���D�9S*�:LDx��2&��c\
 ы���35b-��`�iA��l��F�Y�:��}P�ܧw�G���ge����y���0\��7\EG��e�*�CP�罟��N�<��z�k�uOLӝg�a�P	�+��;�r�xE{�}�F>�xQ����$C��%?��l�g�Li��X���)w♴`�ܩT��/F�)�@�<�����ש y��w����ea�a~����
(����Nb*���v)\�~E/	H�ŭz��?�Ԡ���^��}���������^D&7_���>z�-�� ol��8Oy����}-�[�djGY�� �9�M�'�-�~_��Ě^�U�z�}�o����9I�ᾈ&T=
���/7��*��"n�!]-Y���/$v��
ޯ����i�f�ݐr�^��!t��<��T���2�j^oQ_����u��߮]}'$�w}���j�\�@+n�7��$�VM��'2�!~@6R1��Ȍ�r��b=���f��J��ә#�$�K�-4ݒ(ޗ�}l��؇4�o@Y����߷ �����A �Q2�>��#e�[G~O���<R��!��n��*�케�$p���W_�2��zƌb躪Dj�1������]Z��G�J�eX8͕��U�Ž���M�a�ཡ� �p"�i�^Rm<!�T�S^^%g>qs6(�U�K�8�ӡ
A�~���^�p���o�I+�A�
D����8?EDM�d�"Ԗ&�V�Ӯ�I��a}����-L �M�������f$qx����):��"Fف��j����o�7���K����#EOJz�sC1����q�P]|�$�l-�bB�����#�gX�%d{X���m,��~cw#(^)謱�nMl>�@���yT�S�H"\�ˏz�S�VÇ��KaX�*�t��`䮘_B���>�X�Ȕ�ں�~0��t>.�
mj�6͎+��B� 6��n���bf	�Wkj��L��pZ���&�[�u���*���p�m3m:�-���q�D.�d6�;]W}'}�ϥ�Q�)E�۬X�j�>^�G��G˘�p�@�+�ڬ���(����ΰ8:O�J���ĖL�y�JC��N�!�T��xQ���u���[l�A��O�C�%j�<�=����B(�R��l7�
���`�uf���\ bH8L��������I�r-Mȉ�*RPw���]��:��~\\t���/�^��zD��ފ�e��0��-*����۟>����9z/^��!~N��i�E6�����'�S�U��=�z���{|�p%����U�OMvU@	[���!�$���Q��]�[�{��biU������+�`�)���k�v�7��u_ؽk>Q��~�%_*yl|��a�ca����TG�577}�����-h��k�+���Q�jq?VY5ഝ����3`+�d*,y���,�[y��nN<��J]D��)�U_���� �~`�NU&�s՚�F@�z���������qS�� o�e��yJ[�*Jo��5fgO=��H*"CwR���� =^L�c����	6�Lxu� ��|��R1�b��'B<k���M��&����)����	�	"PO��~ rPγ�nO%h���VI�okq@E�g�ԟ��U`��*���L�xp��
�"i���HiA�a�Z"�ئ�ę���O�cZ��cgp��h��Ls��LT�R�2��vnI_���ǈ�܏{�� O�ߨ���\����o�ꘝ>���.��8��Rw8sJ��kj.u�5�*/��\_a˂_�=�?o��$�YC���w��lC�B��R{8�[�\�K���E�*�w���7 /��U3ơ&����0x]3�e�,C*۵ek�B��X&Ǻ/2��c���![Ҙ�3@-+zاK�-�_�#�~��
�/�i��73������gp\ԙ#��:��yb����(,�
j�L���y����%�@	��@��ˎ���2��}��.���?�j�j�˸
�8.�ߙ�ژT�/�ߘ�<P�������ŻN��	�-A�t�}�<��i>��tP�L���Y�ʾ~�2.�7�{��
�E0�V=��=Ӫ���/#�b�t�K3�1���N��?`@����z�D���$Ѱc���� ������c=�Ы����׏<������<��Z���c�;�2��!���� �u�Z#�ef5/W�`�m�'M�;�#bU���2��p��ѥD#�`/w�����~�ꈘ�>K=O�ݷ&m<�j���u��n~�����\�zt mp|���`"����1}�D�+2�/�Z��l_X=%^l�Lv]�&�}Ï*\aFj��ǎx&m��0�@�Y�Ws������&A�>�1�Ui/qs��Wb��UQ�s9-����}��Qf@�:��B����lA���2��͌�y��m�5;�z�޷�.��������ahm�y?#W������!�3�����T	�q�ά����i�Lu�|�h�3�c���U���M�?O��̔	{
}C�zu�s��ۂ����Mm!}(
�������uD?����\�����s�˙��{�,���:�XШ�}g��@APVN0�����մ�E�����<��R��GV

R�V~l�ϱ?�^���O)����l�<��:�����uKĵ�'��`�$��dr)�.��FID]�zP���LНC��/�\���"(gv�ٮ�f�o�S��A�:]V��;TrkZ�~��A�@mq�@���i������m�Ⱦ��yfMN�{S�U�Zd����V�%��`^���Z�Ic'w�����<,��^L���9Lb��쎑����(&�U@��e�io�!]n�ȱ6�(Gw��X�!b�)ڦ�xTTۨB����K��l\�/Z�o�q�nW� �l������&�,>����2��U�(�M)���?��{��xY>Gt?�̠%x*<����,�(J�R��+��oL���+Ø��c��wo�|,p(3Y��y3S¹d캣�=+��1����D�_��+�W��� 	����8��$bhF�v���aoj�_���y�I��ҕQ�X?f����;� ��R׶��������'�4�	o��6Kܻ�q�\���_��	a�k��6
��a�ʳ
��v��!��k7XD�2�y��P�İ.}4H�\�&��ˏQ�(֔89U�~-sM����M�`�x���Eu�L c{l��Qg�)�v��?!<'�)���*R�q�� �dwIp~�Pn���X�%�8�e�-�4�4�����&-��h�1�]�� ��t�3�ke�=�.���ϗ�k����m���@M��H�m/1��T!���>��Ie����3����u.Ļ�n-f3�J�:�ʼ7��0���1�8��g��.�h���Ȃ1(��J�ŧ�c��PA�Qǲe'���IƶZ���j�52� A�������xO��L�[� TPM�6����.�Q�e�}��v<�S��
^?vN���������8H$�L+}kbJ�Bf7cX�B�\l�J�3�����ȷ��M�ۯ��T�~P��T�1Y� �zo:V�8���v�~p Cf�;�>Р׏���$���p���jJ�5����I/P�{v,���^??Z�*u� �2բ�j��.�"3F��<s��F�<%���<z
k�8@gnX���XF�X�*�!sZ�퉙0WO�@��_�-�[2O�[�^��=r�+�m5݉y�>�<[�NGm��Z���VOn�+�$�G҅ 4R�VD|Ջ��o��ʄ�H�!�}���x2
$�O]���b�t%��׻�����!S���yB;8��OGϘ�p�Z�97t�h�ŵ>���!�2,����_�i�B.��틳/=Z�(d?�H6f�&�9Z��vo[�hL;2j0���Sb�vS�N�FG��X&��v�C������ e�R���'`�BE�;L��x�7�	r���~A�������F���MJz�Ci���(�'�,�=y��SW�0l����ۓ�RLY|u	�8�Yh���nf[�X�ڦ��
1�
��sUd:����E	��<���<Q1E'eM����h���}O�;)X@\1p�4j���AQ(� �YG��91�z�����Ў�H��7됆�H�:4x�> �ɱ�ڄ<C�տ EP�)� K�s󔸩VZ�[�)�#r���T�pӟw͝�P��Q*�W�
�#��o�����b��]jo!�̬��
��w�)k�G*r$�2��J��ǏQ�`s��!�?����������r�A����;�UA���<ٞq�A�x#��V�n��r�<�͖�mWF�
�L3n&j����
��
���R%���:Ef��J��ÿ�5�O�ɂ�]�q�@qZ^�:FIFW?��u��ILvC��M�߽V��;�#<W����I�N�"�z���})L�d�∃���s`��9�E�X]�C ����ՄDk�T����z���~<����J��Ob
-z�9�K���>S�ٟW!����a�6�<p���P�Ds6.)@Ԧ�٪�p4r�3 /�u�$��ؽGf�t�>�ws)�x�L�fy�A����wF�oѸm���N�F��ɇr�AL̎e�(oW���$��hpB���p��<�H{�ѿ4`�}����.x�?���-�Kѫ�/�m��v݁�?�5�4��Xގ��&L)5zW�`ypD��5*���L��su����BP��R�<x"L �x'��t��t�ٟ��(c:^��l�3[�}��;��uz+���4�$4��d�<�"�j��m�Y*g�{�9���<�(�����!��+�>��|%��8�Lz�j�P~�����&�:����ڋ��ֈh��̑�@1�C��.�I+����,�M"̰qS� }�Rt��U�����/��X}�̭��]�Y����xө3s���R�s��_ؙ=_s{��ʎ{{�����k�ɷ�)5aW�VQn�@ӥK���/M�X^c�Ŏno�j% �����6h&�=�j��j?�V��*�+/��n]r&O'oT�>δ)��5}Գ��2�NW����o�[q������.ϩ����')����M�e�Dt���_W�<�	���?8u��(0��T�I(���ԙ
�!:u�[M1�ߐ-��L�8J�׌rX����O��ob���P8�W�c��B��Y�>�	���7��@Z�������ax����� 7��\�Ce@%I�+�?p E���H�ItcV��U�/-MD4齾3�G[B�t{^ ,4&��A]�:n����y1\��ÌߗT�2K a#��;��hĘ�H��xU3�NR]̀�]�2�_��6m����M7�忸	��n֔��K�^�UC���@bZ}���9끨��J %�qE� ��gpYm�[A�zq�7�v� lۏ��~{�GE�7-���F|���]�������:�X��	+B��uI�e������뛽Y�.�R;�g�|�<Eu������ e0���NdJ���K�,[t�~��Ij�O��*��;�ܷ���g��F~`��8���6G��3:%�?9�l�g?%����{���'���#��ב�SL�M�__��xkd�YFh�]�9n��}i*L:�Nղ����t;���VJ��\�`ݻ�`�D^G�$k}�5?=c�cn�2$w7n��?r�c쯍��JQ鯩��E���Q/�!��%�1rtS��I����\��EL�K��r���\Q1(q�cH]T�פM�c ��|�nU_�*���Q�1Ǟwԧ]V��.sS.㴳�＆�ɞ�p8+��dE�+ O�ʶu����=a�:�i���4�����^3�5����\݃��w��Źz�����m����h�D3K�D����fy7�?EY1�]Ev�9Z����h]&Bp�H�/�QK�HE{��^�\Q3I(����`��f�C�N��ޝ;Zɲ��Dc޶ڼ��Y*|D��@b�4a�l8uى�6��������T�Σ�����ڠfV�f���@�zMm�z�<hs]��o����b�\d?޸?�C�Ό�.�qJ����ͭ�H& \�]�q�T���?�����&�L�s;t�l�?�����m��
�[���۷6cc�=���fhv4��������z�x���|���)KR�$%�%YO�%	!�d�'Df�t(E���c���5�0ʞe�����n0����>�������C3���}]������z�/
I�2@�◭(ݎ�פQ�۽���*�ȿ���f|-��[�V��Wo�R�3I,�I\��J�8�|�5�Wa�Y+�J��]���[�T� &:YRH���`7��n��H[������h<�n1�u��!��&z�}�����,f�?��V�u��C4���)k���J��d�������.����^{��gǪ��6�=����s��G�Ro�H[�ͪ
p�r^��P���r ' ��[/�#��.ژ�s�uc�B���Ǔl�A�up�:�Ԍ� _�m�q�XU�C�Ҏ�(�}���ϩ�����fV�P�I��a�!BUՙ���@���
!��\ۓ�c�o�ܙ��.9m�=��^�D���c�j����� ��&u�w."�W=���&��d�\�f]����G��Y��0.������F?*��Sk��]�wECx�;>>�Ґ�;"1!ٛ����9�+�VD�k�XgZjA�/t���d$����z����j����O�4@�A\�����8�5�Ur����@�@
2l:�*��(D_���:
�I����������j@ ����Q0���X]��I�E%�ox���3�p��8�۠m@<o�bPq͓Rv��Ǉ�[�#�"HlH M<l<������=r]C�rt�����a�L!ߟk{NU�pΌ6<qq1կ�M��I�N��ay����΀RQʧLX��;����2���\��-w)�?��'U�K�?0Rs���C�~�0P��$Di�+��L�Ҿ�TlU�� ���󠫘�P�	�drI�4E�[_��X ���B�qV��w�h�91�^o��l�fS9���S������*��<@+�7����s����ty�̥�� c��Q������ٲ��^ԥ���"N�0�<��xrU��t�}�����7+9��S���C���:�C�EM�v$�(�ٖe*\�)0��Â�hYYY�c������ID�pY�@��*%�m���jӱ�z���u�!.��k�̏w�y7�u���J:C���#��������z����&���a��i��������wUJ�=��mӍJI�gfc+���h���D���$�ښ���c����0�vPo9/{��[�y?cx��!�������L��b�J����vC��������/�������1K�s�į`�qBE��d���i��s&{[4?'ޅ��!Ấ�ib�@�n�.�r�Z�c�Nr0���~�����m��UNPC-m���-�(��L>�M4Ց�G��,Fuj3���<K���͸C��}"�lc�zI�`���T/����Q������L��⥖�۽�$+9G��0��ǾZ�h16�D.=�jϔ�t��K��Ѯ����L6�3Wl��t#��{V�3��!-D9�������(̄�PAa)�����˯ɥ'W;{�dw�.h
|���ht��-oxK��������50PB0��r��>-�?/7b�]�	�h�Ȣ�c�Hv�G�O�ٗ�6���T���q�O�q~f@%=�fLdA��G�	�7K�U,9��̍�׽ �S����6�z���d����6˝�="gc����yLZ���[�}>��#�/V
n�]_i�����h�p���^ �[�%ĉ�/JsH����	JVɰ�s%�{~
��L���=H3�Eή�a2���X]�҈�O��:�z��M�8�X�����y�6dOv�}�h�K]a���� ����M�/�FR���Q�'pu��J��J��uDD��U$-/ծ�7��1s���;�B g��B������!���_���{6��P�v5^ۉ�Px�K,K�8���ؕ�����.�yn'��T��H���_�C���Z����*X�WH(s{�^�֛�֩���̊R��24��<����}�����E�c���;]2������j���p5yX��y��|G���j�0�(W��e)�SF� �tKj���h��7 ��*m�%�C$L?Eo����\RX��g� 6]05卝���5�߷΃�<=��󥫫��(��RW�;��J��B?4��1���K��L��I��!��cL��ǌv�7:d��ʨڛIo���^"�=��)!��{�5@O�p%ۚ����]��T�XI݋ʀ��/WG��IV�+t���[�: �<��F��5ݩ�v�?x�ִ���[cϔL�N1>�E�����x��|� ����S��ҷ�S(��eHQԪ]n��?g�����_$��ٗ�J���|�z�#W,#7��i�O����7&sY�)���ߴ��2o��kl�
�^��b��mպq�Q�S��]�:���/їL�&��
��vO��6ٺ��"���'퓸�����Ih�I����}������{��`���3��w��Xt�pＡ����J�8Y��浦��{/OJj��Z��鈌P��4�.��/������9�Ō	O��2�VP��5r�0�j��|��Gk�9���7g��9E���aD*����1�d��Ȱ<���H����Zީ���m@Eu��+�'S�vڣ�j� �/�ڔ�\Is��@)�t�A��+1������be��=s������+�j�m	H�]<�ut�.�������χr���+̭�Z��H���q{6�8�漣��n���)���V����с�i� Z���z�<ڽ��
�`lѩ��s_�=x�}��*" ��F�OhiZ!u�G�j������\?�\~?�(�$reЖ��)W�'Ⱥg���$�����4و�W6��;j���l�i�N�`M�N��+ks��93�ӹ��I��F�m�s��SF�'T�)�pk�f�$� �R�p�dc�<�t�*D�*#"��i��㼑�E4�N�`o;��	 $Zi��H�0�[z���q����ߚ������9�%1GҸ�밬TI�ҰR9��)쨧,�S��f���f�91>z�yiB��7���9O�w����]u"�/>i�c�G�Ba6Z��d�������.�������e���L��Wh6;G�U`us��g+c��YG��k���ƑS��,TOH;�%�)���e�F$�A�P7�oM�Rk*-���k�����
;��XDA{Z��Zx���3;���EJy�	T�����С��E�*���3��IV��ӡ{��>|�λر���h٭�:�z��Ӫܾ��V�G~�8@<��1ض��U�#K�a�hVK���9G3o��2�b�RW,0�1�B3sd��c$5��Q��@�W�n6�xy]�_��Nox�~d��3w��Ґ��T�����S�>T2#�P6F���{X�B>rH�h{�|����R�R����	8 �]�=k�W�DG#�-�/�>�@OK�E�x^$������I[aw��:�ph�C�	�w���8�Ì��D[���=ȩA����5��[S�2�P�c��-���}bɐ`��dXgSl�5,�aL�+<�(}	a�����x[P���!'��,Ÿ[M?P:��$�-ӂ$s �s���F�(��h'��cƯ�
�mW�= ި�1\�X�?Tk�)JE�u<i���ǌ5_�c9��cհ$��'t�}��>3�"o\TS�^�%�,IR��_�^y����)��s8q��F�/��i1辗:��È"��3[ߛGX�����xU���H������=�=�B�!G�hFҋY�qC�g�j+��S�A�R<C�%6]98�����熘�_�
P�`��o�S�_4;�;N�ũ.?>��-ͷk�����h��Dm��
*���s_����a���:Z:�$Q��Q�����Z�PaDF�>����5`w]0P���XV�U4&���mL.Hx�;~���X\"� bs��>!���a7�1����� E��:�S�6[� �?T�<�����*����[)��#�r��N4���=�D�J����`���4������YY�̡��ry�ķ�&`E>����k��˚���ƿ��I��؟�2��V*���t��Y�i�d��P�b^�L/����'�����f_ʕ���#�弲d�� ���ݪZ���8�_��:i���3F��1�ՙ��z>M񭄢H��L[���+�KoHeQZ�<𓻮x�'O_L%of��N�	n��~[)#��	���Y7
��k���3��T�*��]7����D�*���g��g-?�fl0�<�4�\VF.���]�M��HIp�B�>��Q�m@�'��rgAjd�m��(�,$XW���5C�!�l�>q������2�Ƕ!
��^x��%�?���~��_>�C�����׫������|��|&D��'�j*�e�Le��k��;~��@'�E�0��`�����\�^�1t�_Xaы�@��z�4�Q!��̀��0�ڐ�t:�Q��BE��F���2 �uG|���or%øV����A�5�@��h#LnV��.��1mX��\9K�.Ķ�c:�S?W��TF{
�E�e��O�l.f$�8l��|����"���(u�����l�?���D��Z�3!fݿ�ʘ����H  PR�Q�yώ�N݁7y�2�S��1�ۈ*�"׹��k*]���x�@y�������{��,���]�(r�w����06�>g���F�l�ߎPI����%��(�V�J����$0؜��N�47���Z<ƪ$�f]45d�G���f��sfQ����F�k5ǽ����)��-T��#�5*��7��d�wm�ƗQ׸s��Ŷ��J'�[�A��ɮ�[Wz�\��U���	�Y8f]��"fڲ�#���X���!�2rsZxE��Y�"��"��Iy�Ƃ0oh��Ȧ*柂m�����_K%ړ���!���H��3�}�j�u�o���ző��N�1k����>��Tk��/������M�!�`�ᡎ��!:H�����?.�����=�H��6a{�}� ��O+��̣<�� �#_ͦi�0!
�.<���x�Ʒ�)h/,p%�=��UȜ��]u�c�4����e�����Lu	�||�޿��OӀ���R����&�g�]��o�r4ix��ͥ�{/@Z�5��c����k���g�yz�,���4�plZ7�.aw�>�_ڢ�ɿF��Xmf���(��Y9���n/�l��5�%��ɿ�a�G���)��)�[{}M��M�Dwm7����[�l]LYg
|�{m�|�_7�����BEqv�-��-2���'{���2h�E6І��r��� N���Ǵ���/j�(~]faϭ�
��o<��.���Y���#�Z���͌,1ԑ�V���7�N
D5��F�z��$��L�d�����)��Έ���Ԑ`�lU�F��9���Gzt�\¶��Q�~�akf�U9��b)oKB��>�M��b��-�O{�V����P�%����L�C��c�d����iP:��iC�§��/v�>T���~lk_�����������B�y�衱�y��{e`��k.��=�#�����AN���|C�hL�����W��M�҂��IY��m����#���'OQ_���W���|��'���0��yHN}8I� _ ���J3���͸`�] �����������9��`K	���O��T����M3R���Rٲoǟ�sp+�?28d!$Ӓ�ٝ��(=v��\���~��%�36Ç��Gu�X}�3��7�B:�Z�`H��W�FPiq@�2)Vzi�����>�]v+��3��}oTˮT���4%F���ݧpdn��G���~��X��Q �bMw���
��TLT��}N+�}��VИ���IUv�\���}_F��0�z_W�D��������t�bQ�{	XE��@'-�o\�a�лGy�UJskP����=F�����+�y�#����L�'}�(꩹�Rv��|y���0�0'\.]I%[H\����sD�D_��X�ke��T�I܂�(0E�
,�K��|]fW�A�U)8]���4����^�oQ.)��_3$�E?�7yY !6 Q�  �2x���7\���t�J���hz�jB��\5� �hh�������F��]�2t<��bJ{ߊ��p���Btѹ>\�������̒�|�v�.^7���b0��	����#�s�V��37:/x��$�d�NH���T�@�^�"%U	��X�WK���XcF����$��wDF��#y����Қ�%�ز�I���1C��|hV�h�쫬-���>�tN.��	��G���z�D�ҫ����q�d�]��ޓ�k�[r��B{�t��P$R��W[:NT�d�	b�W�l�N��5���{�a�#�|Ek�D��_]U�n�7�::Nn*E�a��(Tw�9n�H�σ��˿]�1�K��,p�..�ݨ��_;a�`>�k����YS�Hmf�z��V`R��x�L�2�W8ǿ �{aȷP�
Tԙ4ϩ*ϸ����ҽ	LzF	�cs�=8>0����؟�N�Z�ȧ,�Z:�s6��̻Y���I�%�I(�9Q�Y�������[�8~p�Wܓ�Mh�s^�kX�QE��`��z~��w���]u-C|j4ȩ���*��qc��F Ή���p
�.���V��d� /{��Y�f��e�傜����YY9�b&p�-X����fg9��ղ|�S��Q���G���?8������j��~G�b��lw]h�a��A�ä[�׮��z�c�Q���κ�Q�hC�ʗ$,=�sA�+�f�������Ok1I '�݋}�����a�f�B��U�j�6B�����A�X��-OMY4�:��3������;�yٍv�<��KPh��)�
@��(��q_숄��k���mX��ސ��I>]�o4k��4iWK��!j1��U�X;�gL���j���&S'�Ȩ�����-��ʃ���$�����h���3��$�0��e~��
���m�Lt{��;�]�g���4�>���y\Ǟ(�jAb(S쳂�&C�)?[aP'�M2�y�iwV	�5灴��Z\qvG��q��������`o�p�fP��aft�E��s)Ί;bF>c}'�mX��!�Ht3?5��.�x��B����\B�*|Ԕ?zj,e�KH�\�c �
p�GV�{$����c����;����������BuXJU��pi(������b���=I��D�#�{V9�� (f	b�u�s~�O{��/�Ma([�}W��6�g��$w���^����Р5�j�uޥ�Ī݇���sZjIg_�Ѐ��~ebH�<ƛ?��U�]˃{���,���a�/l>�����H��څ����ޚG6��p��#�M>Q���Gv���!5�@�!�Z�m�7ߋ��Y�r��&������z�s.�q;����!�h?O�F����IQ�*��s�h�B�Zm��9��H��4�!��	�L&[}��0y7��}R���ܵT���9�;�Z�K��9O�t�M��{�쳥�(5y��{�@y;��@�f�h�ĩK��`�5W��'䄼�+�G�]����`?%h7x� dN�]ZfKv�Nc��7ukx��m��uU��^X�Uǁ��ȇ*���94A?j���+�+?;m��-<��}v��":�sB~����3`C��"^b&�	6_�\޴�PGzO�@,\wJ�:�,3PN�zZ�DdU-��q�%&�߾:�% �m��|0���QD�ۯ{e>��:��A�/�*�DÊq	k��
w�U�ǝ~����u '��}l?��F�y�Qh���w��(�9�E/&�*:��e���`R������FfB��黙�F�,7�`i�wJ��CC���t57�ӽӼt�\�Up���C[D�J+-$�oA��Z�B��������2�SO5��Rd�Gi�B�y5d��AB��|�5���/������c_�v��z-�y���o����}5�-!�s��������� �ޣ�P��a�+�����ot��k�>ʽ�h��Y�} �WO�*�C}ǖ�rG��_J�Q��6���n6��dH���2���Y���+r�X�+leCW-!VF���F���X�+��]��a �$�D����q����v��*2�Y���M���ҌM5G�����Ի���N�P2�1fIe���q�G,�D���|�ĥ��Gr��k��'�}Qꩀ��m�:�5]]t?Q,�a�4_gCx���wp�mB�5��~\�V*;f;q����PkB����͠��~�^�P9?�2=��+�~�A��tŚ���T�*��x�AI���;����~3�#��*�lҤ6�2����ir�,b�l��aT]A̡��6/�#,/�;���afiV��ˏ�h[��	��_�����uξ'v��<"���&EF`��h�t�X��ȟ4y���գFc����������u\�>r��q���|d6�	�n�Y��L���K+�G-�huU�+���L�䚂F�=`@1y)��}�Ku�N�
�<�$��5��?��q�*A���]	�^w��� )O�(�yVfk6��������;��D^?JCp*ߛg�"�c����*h
�.\EMb�>���."�
�}�v�����ǅ|1�LDf���%�`���~��g����!���O����]#�|���������R�G��,L� ��dCQ� ���-B�?�3�bJ;=E��rȷ5y<��R_��XI�{�ǳ�ɞ�EW-5l�����A?b��+��[:�j~ .s�P�o�v�a��m!�?�\�^/Ᲊ�Lyc��qGD�KЩ垫a{�Q�x�.�i�1����+���
���<��~���'�'��\N�Ʌ�]���u�����۽6}�3�=��U! ���﬜a���A�t5��{�m��l;y)u3S�RL �lYl�R�F���*=E���>��X�*���^��K�q�b��#(0:'�He��7�J2��eUWaom�FH�m�nܲ$o'��{�1HS�D\�h����3�!Ĺ� �Ѕ��٫P�!� l�ʢc�������g�0�Pz���5dm>���NF�j�!4W��Y�g��3[AP��G���P���a���_���}c��4Q	q.Kjd�C����G0�*�ֆ5�|$:�[��k�t��*<?b�>�֋3����"u�Y:V��!0����=��1���~8��Yf�� HC�����]�BT,��yG�p���"��x���7�W�(#t���݁#P�����(Ё��
��7��y�i���W��A��029��"�N]��L�d���e,�e��T�����~�;���������b(ޓ�
�f�Y�F�0��n�I��xEA��?|�Ȥ�E��>5(�k���[xiDJ֛�y��r^�J��f�˚�ԑ`����/���&1cv���=	��T����~Mr�_�"��7U����Ǎ�[S���kå4f,BZ�s⇛j���?�Lص��ۦ����>�v��f�bI��f�o����<!��F�i�zL���3�c"b�LH/a������u��Ь�n^�+z�Q	��w�	�X����u�5����,�O�#���knU}��sR���� ���h�T�&ybm/BMJ�r-�V���'#H���9*�X~�(�|Zjp�6na���� Q�n�)��"�j9%���~k+y>W�H
���)�5,We���'�eq�9�����8EV���c�\32
6*�FҞ;��C���;�L�����R�w_%�%�qy}�v��?�)4��(�"�WB�
�S=���;B*�fe��Ǣ��q�F �����y�f�4���x���$�M�o��.�@R��#���IRV��3պj��0�7YC���p���`�/=��	�#���PFy��_7،�N4zg�X�2���}j����nm�'��d�-���g� ��z�y�$�m^h�Ӯg�&�8�zW-�sy�D�[���ﰯ�ӍlѲY��k�?z�MC���͈䛐�d��gs^���URG���S̢�*������U��q~���-�=�<��\�"�@�rnl���:�q�� �T��N@Y�ƣ��5V<��O�&ł�yJ�6��f��Y(�2ǳl�F03k��2���.�5F��<��Ai��J��;��ÅRQ�3e�t��<j�F	�%�
ɢN�Eʬ�S��ٛ�wD:�]c�n��R��K\#�a�AA�
�g�;�n�|lG7���|N�˩ 9���!}�Z�@�?�,k[��i���	�� N��`}��5Oh��Z5�r�"�+L��|t���A\٩�#��=b�y�@Za�"�JG�Q��J�O��g#�z64�`b�מ+e��Rp$ɸVձ�_��1��E��
���T�jKf�Rz�Gݙޫ��
�!g��^�� :d��8�S�0J���ѻ�eԕ���;x~�Lb�%��Zv�Ղ2�!޶�r߾��R�y����0����S������s�*��Nt��Fô ��0����I�d
!�Af���J�p����w�}De��u� �>�B��n���C���rj��0P����u���~	�V�i�� wvT���'��D8�a�i[��Z��2�f��د�,�]��J��h}����i�=���k�4�u��^zIJc	-�ۧ?���Je��� ��?��u,6��/���p��k�䨨��9��_�0lR�T."���wy)T D����ًxC�#����^c6�F��5�wh80ŋ�(gm�&�6ܡ֌�F��O��i�+�Fu�|��c_Y�.�?j���W e_G���U��%��0U�������'�=��Q!��:��0к/p����h`�<)H�t�Ó��o���8^�=�ZԚ�6�w>j"���;`��%'�MjBSP;����G]Ea't��"X�U@a���Ӫ�C"�RrD�q��U@�:���~j_2/ $ ƥ��c4ߗ�yo����y
f�R~O:_�]�5TK��<˰4i�c���&,)n�f����m��~�ߜq�us:�z\�Q�Z)��t߻s
��`����fڂ� ��4|�8�㑵;�T%P�G§=d�00�����i��[���=��u͋��Au��� ��½�^Y{[��Ǧ�}�K���]�����6&�m��jI(U ��#~"�O�h��o���?E�o(ik���e]f8�*"'�2���q͸���m@�L�8q��`�#��XB����'R�K��h����q��Gػ^���	r�tU��[t���В=y��'G���y� �����u�R:9��u__-�r14_@�w�0;�v,{�� ��W�'�����g�r�7�T���,�-ͷ�YZ���k���m���ө>7jB����5[9]C���I~���ݡ��#�{��n�e��w���8��I_���c9�^ze��"3b�Fo��X���Ы�Ko�[�>��l���Ag��z�}揺�o	����̓z���J�<L0�agC�h����1{�AN��A�~��g�y��E���e�C޿�� >�Hn3�WE^��d����i6ŗ�<��/��Bе�А��4�̤��]m�M���X�. +t`��y�Qa՛ԏ�~� Fn?<i�2��#���������\{$�lc �Yd�Ճ^`@aq�����p�.k5��?]���ޯ9�Zq4'"�KC,���L����Hw+�Qz걐�L!��OŰ�V�Pnv�sO���ZS�T*9�^s�Ї�Z�K5l\�~\C�� �4|�������(:�p�o����po .z����	B3��6G*w����oʬ��)=��r�Q�~�� BG$:J�a������п�t��l����˵�[����Ea���Y��-
��+1�r;��m�@N�8Si�_c�Aƃ�Q�(CMq�4":��z�#��2��ǩ�����#�0Z�eK�M�.�09$i���|6�ǯ*veVա��O�$r2��r�G2O���t�?T����k�lcbD�. y{	`�p���w���ۿ �,_�L�7���x&�v�e�ʷ���z���L�~��Tg}�pp�c+�P�D<Ŗ*�!�O��$�fg=Ůq� �$d�-�L�UP�ap3l�1y0��R��pBduv$)���5�C��i�/L�`��)UَZ#��_����j3ñ�",��|�W���`t0��]u���)�g��N `�\|T-G
���P�����cu�cjl��|���m��&һ}�0/R���:�M�|�\�]�����z��%@xw��f�i��t�aq����=}Q7p?������_����y ��jȯ���l��v5���5��sKbb!���a&���L��0���-�u�BX�I0��G�"�/	0G��H�(~��z�/��^׈��H|�`�2&��-D��<���c���KHBE�>�i|�r磛k�D�����,~s�
JOBE�`�lա��ѩj���*�r�?������;���3yc	2e9��A�lLZ��1���L$��")�Bc�o69��~v���hU��yYm����� ���pEg�Oa{Db��	D]+�&a�"�p�Cα����GJ�߁��.T��<����Ț�n��SͱO�V#�(q_�{�u'b��߲��AN�p׿'�:D%��G�f ? nM��R{sd�&�J�s@I��5���k��`�q�L|�pn�Pk�Q%�eY>��0L	��X�~��:���{�E�B�K�lt���s{|�r��<C�j��� $�)ʁ):�U�~{+!zb�`�r���@���{��A���+�V*�@��ܟ����>�}qZ��F�R�|
�f��j����a��{�Re��5�6�LE����|�E�a�Ǌ�w����'}��D��~Z��4�=n�x��.�о��{ˀ	�}�ђ<�<��m��\��l���S�	L c�*[�������: t�7K)g�H���F��Q��A��h��Did���Ah� ��@g�F�DѸ�5uJ�N/9Ы��Y����FO�#7�#���<5�����wf�O0�9�2������}��iԂ�f�r��2-��j�ɣv�}�x��;�"l�R3���V�r����/��6"@����G˯n��%+�j�&�x��W�-u1��x[�]Wyx��@�Ia�iP�Y���>����������j⟬*ƚ�9�s{���D�g�u^hĴAUh��t��dj��&�����`��;��t]it�������FP�pfmy�~Њ� ���J|	e<X<;��F����֕@Y�y�F��r���hϲK܍�A�݁�N�\g�H���S[�2�� ���&��@����e`�������� oy��AC������"B��*�_+>Jq��_=��u��l��sGBZwT��%8k�X/��RSznа�������0�KAT�S&�xtw4�A���;��������}����1��o��Ε:���S��i�����a�c	����0�8�9(���R`�,��z5H��W���պ�p]������5�Q�߲A �K�F�[��t�Z��%T���JU��~'�n��Nz���h�@Q*<;A���B�U��
�ː��e��{!�*����N`�U^Z-xܡ9\�jr|D�2	��$[���@��{p�KC����2z3��ظ��<=�*�u��a���X^�OE�����ᣅ�ː�ǟ�~�H覙��s�2�-)���YN�������9�o��B�!M��{��W���{�5�9����Q�/��M=���N�o!fJ�#r��Q�IAAD&i��R��Qi_ ���<��)g���r���㹱�.A��3��k�� ��kW���6v�-] ؚ<���}�W^hI�+֧����]�d�����
n��G'1HQ�i�*0Ob�I�ӡ���@7���{�%�O�\@1��2=fF8�&��d����}�E왜�jL������#~�oߟBd�w��G^MB�n�(��5�J1���HL-���EqA�B��I^���K�{�$ʤ�(Y�ğ���n�e���8ㆬ
�Q"Y��������^ڃڊV��Z�����^(���i����Z���=ג��2�����
�#��H\���_��d�T40�C�	��V�%!8gD���5~koY����$��ˀ�e��e�y-��Eh��y(��!ɮ�a}5{6'5*n8�M\���Sޛ���I@��;�NZi3	��[���:�Rשչ+��t]R~y�L�3X�͉���0?I��X���;��%L6�zo��F����y<r����2��3�|������j�*w����c��B6����$�4�eu��Ũ��!A�x��9'��GUN��m��_XK�-ޜ62IЋY�-s-�{{�.Q�H��:�0	���O�\_��M�l'?�V1pe��;G.U����l����v J���R_���!��k��Y�ި޶pQ詩:߷��1/��	t�4�Iw��:f���{�^��m3��hS_���-���*���Hp03�X͓�:�C�w��;���N�x�B���xa�������vVӪ�����_r�\Tg��Դ�,f���V��/�۵�M�n�x79g"xpk���[DB�Ϯ[�������:��~wD|���ծ�ׂKg��)E�=�_7����sԳ�H�����8�o�@Ѫ|vb�S�Y�i����,����<�ÇǢ���Y�'�.q�ah�9Y^E�!���>���{5vغ�]���ͬ�}�k�=/M��Ň�g��x,7,&k���&̮(��zk�R��n���sU��ͳe.o���<���	�~��⪗�i����,f�����v�L�	��#���<+���H���\sf���X4��KG��	C
�/U��o9�г��e;�%�����1AucC��3���/z�)4%�-a�M)˔?�� Rm����血q��fy��[��J���۟f�P��Z`mZ�8Y.t��vc_��Ib_�R]gɭ-yC]ͽ�Gڊ�����s*�_��KXaM���k�L�ه��6Q��ܬ���NRae�C�Pu?�8�#o��d��ϼ�ڂ��˭�Ƽ�Vd0��w�|�P�d��Z�L`�U^�r�i�X��	�S��~ARy��I�ƍ���J�ک>�s�H!h��kƹ��{UIj_��>T�g@z�Q��G�rN�Io[���r}#����z�����J�^uO�'�*G��GW�f�{Ͳu�U�����b�����e�GQ2�=��.>��:J� �x�H�����wF>!�Yv%�Yp�uH8����/��=��9��K��-U�ٿ}�w´�vbX� �O�����q.�o�v��W�o_��mN�Ζ�t�ԄT !űܓJg�W�+���F)u0��S���L��\���{�H�����=�oMc'��4�N�����	!C;B�t��R��t�HncM���,�����7as�b_�J���l�J�����	@����.�	�3��d#��C��[ZOD��6�$�f� qЋ%7T�r�D�[~7�����^฀�L�Jy���b6V�5��`�w�w����Z�I,��⣀X�G2O	"�J��L�J�t�8J� "!��������������:��`U�Y�D7J�����ݿ5��KUWI�̱Q���sU_�1P��0wK�!���=���e��C��m>u�D�J�����^�Ϣ�|a-�������ؤ�U��ٳ��"��[c�8�r�C�]U�
�z̬>a��o����Ć�cy�g?�kr�r��'��~��p� ��b�����-���8Y��;������-l�L�wS/q�>}^� v���� \1@�czο'%�ױ�����P�-{���qA9HާR�DN�g���OY�1u��o�9?&�a���П<j�@�rk_KWYj~/��_��;t��*�)��7�'"'������6�ߚ�5�v��Pzk���L�ɭQ�B�4�.6L�w�4?��~~������Z����g��+h�5I�=jn���(�֎�����6���'�O�>�T��3y)[m	K��;ԕe��f�&����Cs��b'k�^8����N��S(�,t���p*�c�w�n�)� ��I*�kO�����'1?2_��p���c@=���~����P���h]�z��7k̕��,��AP`y�S��z�\�u@T�n�/!
�&�ylXW�4�
](O��k+���G=/hv�BBkX,
MJ�Y�^��%��9���6�|�fN+���u�� ��|f�U]���o'F���B[��Sz�Ϭ���z��N�����s7H<Y�s����@>��B�/Q�:M8l ������7Z/��F,�����V��#�3�%���3��h ���^Dܤ����Z�~��I�hP2$WV�����Љ$�~�֡��ّ��cl�ky��@}|�V�=�/�U2u]���>�"(S��56�ڧ�͗ҶU��S_�a�SR�|4_���D��Wm@g��Q���AD)����!Dk�k1�����gD>��ń jWN�����iG���8+q� �De�*���y�� #�!H��+����-KjV�d���r*�X1������Ԣ$V��L�|��qNeV9���2|�z|���HU�-�<䀛�g%�zQ}����dTd��;.+e2��Ig���;�Q��l�)L[4��ۑ��*��~�A �<5��*�0m���-�N����%�ԣ�|�s����w�^Yn�\x���;� ��,��'����n�G�x�aƧ�g�r*��A�1��;�Eԏt�������)�"N���%\�B<}�\oyo^~��ڸPg&ǋ*�jb|�N���R�����A� TZ��a⊭���ۮ[;���D�U�S�-��+��uET(~v��t��-�x�l��kؽ����&��N���<@J�4Y ��?�	Z#u~U�O��k2�)����7<S���k׈�KIquȧ>�if�{�b�%A�N<%=�ґբ��<]���} G��E3�P�Ͼ,x����:]�W���?��h*�w���K�Ebm��arx�>}A݇��u|��A��4�ؾ�Fr���{c���cv�(<���K;O�_vy[�g�F*S�:��nJ8��
W;qN����5m��������j���@+�.[o����z�)���p�G�2���3L��]]B���;^�������P�q���"$�w�"co��0�~P���! 잳�l���7�>���%�pu��}���׹88x&��t��P�� P��q���,�����^���	J��A�i�נ���s�i����E�j�55���[D�^!��MA�sȻ��Aد�ә��;���f��1���_*r#�s�Ҍ��l��i�@�*r��{ԴM�	\�3��dOผ�� �v�i�GV�Z46D�:n�ZLs��Q1H���V��c��y�a%����/��᠑Չ�Ԛ���b����W�(?�z��R�e$�^Ǻ�@ft��Es:�B�!h�!&�{:��Y�V��n���a��!�;t}����5�������Rj���� 8��
��i����M�����S�U����@@���[w�uj��&W��u���E{��~p�n�`�������:��ײiϪ�� r
eIEb���y��: r��{�E���82sE0��8&@�J��(H�aT@��@���q�$ �b���t�A����6�dhr��9U����_��/��Z�.ƪ:g�����g�*��16��#�>B�ƭ4O](�D��y*�W�s�Q��Es鄉�:W�?Ij�W����������l|��#OU䢸���� 5N�Ӥ��Mx�!M n
����/&&>U�F?�Y�8�>�	��5>�Hf��v-t���Cv��u�Dɳ���>z���'z������L�Q
�D.��j������M��hc�����%PN�1��I>���^�׊q+O����!��|��Z��dX4����� �Z����(�N��ڬQ�����vv�	�j�A�ϡ�fU���eUA�~''oA�.�$u�fs�ʇ�R^/-F>�����Z���A_Y8C{F��~0���.�^X���@R�Hq��H�C��&��7�[����(˗�i��� �j�?P)��ZCQƞ��4�F"�͌��)��1�_R�ߢ9/��ާj��C���e�Å8&�������G95@� B�I�8��4Lw��|� ߆�K{}!��c/���A��-���N˧�xl�|>e���U�둺@���	����.\8���֧�t�g��`��kLl|��8���A�����&�Z�m��q�#7��E�86�н�����PY����>:o� V|�&��1�c[�����|�mBڗX��:m}yױ��HȒ=� Ś�q�}Q��uh�x�xg5tv�Ә�9/���ve��VQ$&n���8�X�n�?���qA�6�+(7��6���2�Kq\:L��1�����tn��.�$G�����{��)�/���F�MT�-�����E�s���pB�^y�,}
�g�o�̺,|������X�N�;����]�ƛ�HJ�7�ThtMAr�n/���j~�~4����P(����(�t�p%r�vH�@>��~���j���Z�=���:�͔�A�r8�H�@�M�����9t��������?A:o��)��ǫ����zty�u"ȴ����)k)c�S=�HsG����U�Li�N�����Ȭ�e�B�dz��5���ª�w��ɚv7P*��G'-�*�� ٧����n��c��oe������4��+��<���s��*�lu�	M.u7K
�zϹ��k�d��x+I�.���bD ����&�Џs�0e�u��N���}�KA$s�x�	s �v�k�(��d4�&sG��u6/>q?n���:��v�>0��� �����Xؗ�M��~̧�k�ae�b# ��_�����P^2�R�h"��l���S�ڦ+�=�O��}m���?N� �-�vay�*�����-yF���!|��#Ӑ�_�����<NG}���AX����9����C�&A� �Wޟ�(��:7ydw`�Q���RՕ�gzz�\}�|iq� �����$��@z��\�r�U�#ਝ�o�������vY�G�~R���@i��;s�별��8��Ey�]����/V�|o��]�$�����+®~㠲6�j�w)����{ޔ(#�0��s����d�����j��|��N�/�nϋ�W��ԓ&��j��WN�� �Y��Křƛ ���jεq����	�╫�"h���%,(=�0iw�Ջ�H�w��#�������p�����g���C�U�]�ۖ��{�QU�j}=�r D����Y6�9է�Sչ��%_J��̏ �	�%�,x(����[H:ICtS�&��.�y�[��s��_�207��W��S��f�Hbu�.�OD��Cn�#�* �����^���R��Rl^�U��$�P�{.i���W�#
R����1UP*�<K�{46Jy-{�����"�����zQ�~k^��O�Q"MZ؁� 5������;���:*(/��C��k��(Q�g����MoJ}gG���S�}%L����& h��AR_���6�__�vr�RP*,n;�s�O��MM��9s�> �ȇ��������W}d,"�#��Tlr��]�ڰȿ �ʾ�N��.�e��N�$�?B�?zT%[P���T{��K,�7;~K���q��-�������������'���ؓ�ҷl�������h������cN;NןY���iX,��o���^�s�JYӣ���f��n$q�Qy_%�ڽ�t(jjEU�%o��u�m8��\]�4�ƍIe�76_�n��6Vx��Im��9|�[�b��3�S�[��W�,��p����A$Ҥy�Ło���K��`�X _L�rX���t�h1�����7�8Y]���&�~>�섋'B�]�k�Ȥ�Ak�M��i*H(B��*�1�e�!I��7���bV?�Oۓ6�^h�uF{Bq����	�U�N E����N��)p�6]�����n>�E'�8��S���!���>���۞[��I��EWE�"��Yx��Nۮ�>d�9FuG�ĵ��"���yu��K<4<��%���g�K����V�Y��S��J?��lEsI��v���'uS���Y���Vm�G򷄽�sm>[@9���ѓ�9|���GWzT��)�85S�͈l���D�����:��,�r��'��%hv~�n�Y��4l���Nhp���\�l�Y�� �'� _8�#'�Z�/�#���ا��9��[�p�E��v/FG�7��>fe˕\OJ���ߟG�xNMJ��e%1ڃ`'R&.�S�`�B��.�Q������-?���i�w�oD���?@
�0�x>ٙ5ݏ4�(o�m�{MB<�:�v�{�κ	��V��Y)��k<����n��o�^�K�B$���&QFs�u7��i.����ȁ��吢�6�!��$6j�i��،QX�X<:�� ����y��l�~��gAα��!�-��_����z+l��m �B�?B�*��Mg�n�:ru�˄��n��]�>^	N�>�f�����+��uҙ8_�''�zW����&�]l���nu��Ǔp����;�ޭ�F�|ҝ�wϪ��/�m���C��L���7���Y)s���'�YI�E���0������l|�!2��:���?{��q��sk�r($�ԇ��48�~uJѕ��#�p~��T�C��l��;͢���z!6^G��9��҇�:���u^H'I�H滤�J��s����$7.x�:?���kI���y%�9Зڱ6zQhf7�.���L��F/���/`FjQo����&�Dy[�f�_I�O�)�]ob��߀����F�6N���]o+7{�������,���g32���e���/f2�"$12���yO���=	�p���U�Z�riv8=���2i�2-��[$~�߱���]��p��BFQ��rH� S̦ӓ���	GA��壟�k���d��- rg�p`WZ�DMsE�#�*����f�e�ꕽ
ܥWƱd�T���)1�(����7T$L�����Nn���|d_��z��z�����v���q�1��NQz��B���k�B��]���G6�8��C�J�A�{I�y=`k�S�A��B� ��w�]�?��/��0Eo��>��e��0��c���Ŕ: �;+��$��o������O4E�먼=O�6mH��<��%������%+���0@_M�	'��M�;��?�I��p�$ǧ6�F�	� i�]Œ��UQj8G��с��y@�#֖V�����z4�P�y
t�g@���q���!�+�S�N��y���SB�̂i����]��2�W&��خ��u{%o��x����;E��ԣ���R�O���J|[�@��P���Y�q�Z��-��d�C�ss�u�-�Ps�L��.A�Z8\��g��Kb-�^fj3�,�31��L3��bq�z5�_q>�t'��3 ������,X�@&[�Y}�^�Z���.�7*ڡ�aa٘?��&��UVeFa�T�.Hfm5W2oI�����3'#�_��LB�\�d��rҭy�6�4��{pN��C���{d�_�G`H�X~m_&A���2Ǖ�fq�3)���,�/��.�u��	����.]��ܩ��+�u��՟Q�˷T|Q*��`��(�&�������(����`���9��{�F����Z��X��<�����=���R �u������y�*��:$)	�o�Q�R	�U�����he*\����>�Q���c;E(ݥ$�4)�q�{L!gŁ�͛	�E�w��D83x����h,,��/i:�A�@�w"�]�u]�ׅ���63����|ݾG�,������欌����B�A�]���i奡��^�A_������3���ѫe�7��<(@����	�9�Q@�M"F��܀[*=F]J՟���I��׮a�1N�%-:��T�䖿p@�#6�v�~z��0P���߯��G��f��~�"e0�qFSO�0�Pl��ˤ�Ԫ��`$�� �J��S?􍣀�$W��W���T:?O�É[Օ��D���m�!}�-��ֿ�[��B��2#�9��>�g� �n.p�(g��<�'����B���0o�%K[��a^��2�Sv[���a���[ ���Y��ֳҗ���MuB{�Sq.y�Z�' ������:���Z��J<§+O�AUZ����Q8i͌����'p�wO�_���~,3�N����@��a��%$��/�vP��[��u+O��i
=��r��ڧ���D�r�mA��#�-�B���d-���*��S� ������,�2���L�7�%�����S̩���C�N Q{!�̯���T�e��7�~�N��p]�ج%E��I�pڀ�jG2�����*$��]I ��$��E v1u�<®��;�\_�E2lC
��vg��\C��K�;o#pY��g����g�k�J��9X�j3��� E�\w���g�*�z]8$��"�bg ��o$)�Lʐ���}�AI<�i
w�$>Y�ʰ��}� ��:��?:|�=�ϝIN�ݏ�D��v]k&A�d8E>�����|I�͋��K<h�v.:�muf%�:�58�ȧY��b�6Ԁ+<du[�x�q2��!��[W��iB�<�� �iݮg�����ӂm��� wn���ɬ%�\D9��-_]O���h�uM�b��� /��Q���_F�$�!.�jZm���w����_qu�K�ɡI
����	�=��,��Q�v���p!��,����"NN�~ѵ<d� ��RAx���=�����k]�ɇ��tt�
+�뷸�;�S=8�L��@n����T���֋��R9�u�#(��M��j���T#� 	^�Oߡ݊�C�=�i#�����#Pa� G,!��}��7��~*���������>�-�b ��:���.j��FeoWQ�j�-��e�"[n�-���Rn:0�Ӎ�^�$B��^�(���6$ܧ�V� ���q�t��b�U�����pokK9@�:*�j�������Vh5���Ay��)��n3�X��^�iZ
7p�J�ƚ\P�A��jƢ�oc��c(���6��9���ihX�V9�|c> �M�z��3e����+��8��Bn#�w&p�����Z�d�yU��,������a�'m&���~4x�RO--�+�N�3�N����E�D�"��j+�D����j\�Bg0l�=5�(g4�ts��+�>��2�Ek[�	�v�ӕ�od�*�L/��i��&�/�f��;�p��$�f���j%�9��
"`�2�duzm�()m%q�4�irr��0lX��{8&��৵@�������ڳn�l�2�����+WϾ��d}S��[BK?��o����Jl��$f)J����嵻{��C1�K+�*3�cZBJ����@�ì�<���89��]C�&]w�4��Z͌��\���cR����E�~f�0���U
�������BPS(�cRj����-/�dBAQ[~���A.���4��*0� b���w��0��n)�_��K��nvjN��%�҆k�>
~��>7k�S����~q=��V4�Ք�;<�����ͼ�f��#��t�#�eU�����g<�T��B3��Lj����aM�' ��6��k����/��o������ �Uc����r>	��P,~�罤�$����G�m�r��
d�$�/I�>�=�����B6�0R)~�����(�ˋ�l�S🖟kY0**hU�
X�%��e�R�(�K�j�>�,ml�P(����8p���4$r���mEd���x캤�Jc�1M?{.�VS�8�(��+ �Ճ�����6Ȋ��K�.G��}��\�|������uP�(Gw����?�v��l�X�ȧPTV���sf�	7Ɉ#z�nŗ���C��n&��ОH$w�]~���P�Dyt�w�C����g�3��t��>f$T3k�9�A��9�<8!R�R�gpf��:��Lu��F��:D���+�����u�����W�&�1&���6C�)6���c�DT	w�By��8�����~Z�z�!&��%#�]���$P��w���ؿ�I��/�� ř9�A���֬��%�Z�{PJ�RJ*�m���*e;*5� 
��U|��P���\�&o$���<��a't'��.׿�����vγ|�p��ˏ][��>n���FҒ�2�z8���_s&6Qޖ���w�we�5���u�"�v4��Ш�Q	��T�v�����p�'�]5i
���q,;S��e����dD��Zy/�6%2!���˼�|o ��:y~$UG�Lo�7�[w(A�	[��ʙ�	�A�dX	�7o�dOqԨa�+����#_��d0��[]�KNÎ	�&�8�39���}�gl2��|���|GM��Ʒ�*�=b���˾���^�%��޺lo{#/�-�$O�2��Q��݆ks<
*D�^�~�O��T&��8ny��c=t���Lv��QH�^�U�f����w%<���<��δZ���<o��w�.��!)ÉR2��B\���݇�SsAƾmf�Hې��~��Oq` �ѯ�ߟ�;�x�!]x�	79\�������d�Ƶ[�Hg���s\��:M��D��g�R�<y#�㰠(|I�e�,m���b]�T�	ŵ��2��.�}�QA2;<�n���_�Ar@u�9��Eƪ-��7��7��Ѱ����%ʿ�i��DK�l*MH�i���"�k�9V~�
;�3B�o���ʖ~��L0��$��L�]sȊqa�/?@&�؜�ޚ�9< �N���GM�7�n��b�$Z�� �4�Sϟ�愘(��*X��aO��?r�PK�EFTJ��������!��O `��
O�qUd�ۍ�W�5�9]�b�LR��G�	ܛ��Q���!h��o,�|-ކ?��@|���5��[E���a�v1���Q��*ʅ�-rی�KC=���@���F,mzE٨xA��ī|���p*�F��6P}㇗�P�_\1���������N$�k�B'���a"w!+�k7o�8T�P���V~7�:�i�U������ЉUO�p�8������t`�o�Í/I�+p[z�C���7���'@��`���cΗ���3Q���D�(�*1ݺ7?"��[���O��p7��U��H��#/Hp ����3�q�<D�|B������w䳦F|U=Yg����̚�\iN)-�b߳dt�4?",~�	x�f��g^t\z<���-��~
�]��vF1�&�B^�|�_����"}��(Jf�qqwo�6��j�,�qH����'��I�.~�-�= �~����Ȧ��D�W�#.0�w;���Ӌ�07q����������)w6�־��($�M�������Y!̰3]H`��R��0�;!՘�N� -��;�LC�i��g��_�Na�2=rF����m���-<�&5�2*D���������;o?L7S�F����p�F~�0Ʌ������h���&��#�!�թ�M�_�o�����1
t�9�,��=R����_�+àl�]P����{שZ��H(e�ȘC�x$�������M�����<� �^��J��_6_j���.b�Q#���۴�y !E<��<Cf���#��{�<�E�p�����ʰf< ͊�˜/�S��HNS�1*�P����R���������d;7D�~�Hƒ�9) �w@��[8��ҧ����r��Mya�nٔ��i]�Br,�'8�<�y�ϓ�֔�;����j���V���`?#9C�ÓmV?�@QA4J�n��	n��Gc�.aw��,D�إn���n���Ƀ�=IW�P
��?�b�$�l`�W�D(g�����E{�p����s�Cۆ�|n��,���e��tDqq G���[��=�0S�뛋b
�y���m(w��R��iE]��|9�i�9�j�:Y��3��Q,If]�t�%�q��T��Ɂ�46�w{��mvK��0��5�0e��:��(�c�f�����Q�$�.�2��E�#�rm&� )+�\]���߿ϴ�W�A�`����*�����^���2ZO3�>h�U��K�������K΢
�T6A#��8�.>�S>�9�ӧ����B	SW���aH*�V@��N�t���X��&�����Cn���{j�C� ����zv����)_m�����n7X�k�3᝻�����L�y�8*8j�x�DW���E�����y�na5*���2�y2�ij���_�f���c�qt���I��6���f���S �Ct���H	f��m��δ��7`%#�e��־��Y���5J奾���)���}�c~�!`�	5N�������EƢ��?��d-�c��OTHUeW��G`���Y�� ���Rq2��<��\���
K��!�֎��i_L�Fk����Rb�|f0�?G$�����ל����E%��@M�$7֕(g 翲��^�G�d�~��BsBWT�H*XB��ڭ̕h��f�5z5% 
� ���7(��zRr� ͅ�v^5A�]=`��� !�grA<�!�'����im d ���@v/�ε!�kg��ȡ�������3H8d��O��ѵ�(	��4�D�s.b�M��
�D�l���,��C�zγ	�����郞'+�	�fL�}s���*�����}p��?,�&����T�w��f1�N n9�:8�N�?w	0�\��W�
P���Eg��@ß��m����Ⅸ9�~,|�+*I�T0Cҁ�<@�Z�����G��a?��fDٯ���ֺ�=��2$�"�$�L�h3Y&��O1j)�{���ֿ/{�!G����1���m2�.�����o�#԰]$ې��/�C��F��{r݌	T�͉W!ַ�'��)��A�1��5l���x�U�L���fp��-/��4�@m��6���܃�2�����'|�x��nm�6�~
S�轗�s�K�@6�lLu�ԏ#�9�  b�yzm	Pa��b�� h��'w�Hf-+I��j>�7�6��R0�T���œE��-BD-9ņ�5*�`-dVW���P3[+}�F-#1�M
@/=є� 6�B�_z\�{'��`�������j�:#`X�d`�%*E�	^�z�)JZ8�
 ��C|�w��fd�G3��R-�� ٽLȗ�	ڇ�����N�:���*d�h�^דe�"_���icV���`�ȔKX����"����(�h�Q�"��xBsY�\��P�~dw�^e��|�SE����,S�n^:����3mm��$+���vzX�E���F�Ov X8�ι ���45��O�e��õ�d3�G(�C�I�:c��m֮!�P��\��5j��M����}��o�=��
d=�9FC���"�]��)�#`B���O���,�8�z�;���;�ȁl�q��D�̲|����[�A ��������:>�������c��JK+Z���� 0�-���Y���Ϭ,� ����,�}�\����}� )֞�}�����������
P.Cy�W�K��k��,��v;Dz��M5��w����E,�"����f�S�|�" ��?���j���w  ,Ew�pml�`~C�]���Ba�L���z˷�g��7R��o���k�t�e�e��ۃ�'�1�o3A�� �H֝�����"��7,��n�[Ѵ=�I�E͙
�"�{U��k��]sr�qS^`�~�r:�>U~��o>iV�Di�+	���LO<���4loe��=�hL�9C���ٞ �\u���?����@��!(���DKuI!���򲪢���@V����Ϳ�௷�� ��w�&�G
GQ]�o��L�{��|�����^w�j�N��[W������bs�"��`^ 5���k�Ji�Z�h� F�?nY7�_�F����ЮV�@���-W@�;Fq��;ia��~j�ϯ4��v �f��jAR���/��a}A(�Q��&���!��|�u�M�
>6{��m5|�du�pd����
1��] ��A���鐏�7���n/lt���|}<�7��O�|�Ŵe(��\���@.�H�Ȕ�L�Yl#q(�.����m�@�Z�2�i�:2j�ζ�>�fBy>#�X����}fT�p��Iv!�Wˇ8�OUz� .��u���$�a��Iݗ�Y������~|� ��oi��fQɧz�Wm��X{U���?������XW-�����^ܳ>�b����=���y@�Mm�	j�i`{)�olEr1���&7/�6��*�2���+�w��}|�Z���@�w��I���F���[�ea%5����pdgi(硐�ζ�F^p�һ H����������O'< \�U�� 1��`�0���#�O���?��Nb�1=0��Uo�E���i#����b�"L*:}q�����`��6�г����8�{|�hw❴��1�8��\A�Z����#��K%MjFAq�L]&C{�}�$�F`8�埳��R�vf���Y��UJ��!s ���p�z��8�1(�E��D�,� </n86�t5�H�~�pfN�|�q/fk(kSdޅ��P�a%��?�e��qf��)D�.��<Q�X>h�X>&c=ٸ��X{:H8/����㏸HKב������������xwD�G �{ԗ3F��ڏ�o�3Kb��o��K�H
�Vב-��K�,����Pi�A&�b��÷��Ϗu<K_�K�q̺��S�l�޻�9OՈ���������4�u���颌��V�x�\`��Hz�wF��uO�������؟�[�d���i4�/>6�惘�Qr��pȪ��r�kౡ�(��kgb���}h'�ߊw��/�M5�h�ixAw]I�u9�Zҝm����D�%ŭo\)S����K���?�t��	����˭��-\Y��9�t���<㿲
+��+n�=o}������er�Y(�T��moV�)��ɠ>4z�]�Ԫ=�H�P1����y,>���n���(��+���x;�Bn5 �*rn�
Z��+u��_`d"�'�,s��C�(���5�~�ɣ����Nem�W�����5m<G���TI�x��=���	تwe�Vp�;S>�֢� +��n�Jp�a<��1�v���0���oN/x���@D;.��8Ca�|ES :eߑ�f�?���(�_zI�Ɇth$Å��t�k2*d�Ζ���'��]Vti��x�G��f��|(qu2�7!LN�cmlhq�,#H^�b�����B��C�48q;���^Fc[��
������ן���&{]5X�O��V9��ڏQ+^7{�J���=%
K�M�x�w۸�x�p��@�o.����4�b �DT�-�'Ʋ�M[�<�u<��dp�PEc�2�%����-�(��������s�{p�����[ ����yY�"�8ye�N����^_���ɻyfI|1 N���7��7��ί4/��0N��p�����~��{}���h�i���Ӱ�k�|L�d��;�F!P�uߋ�p-����zCgI��q[������`y��ȹ�+�3��3���t7���.{��6��
�w��xq��J`V�
h\O��t�ֹ�0��S��]�Xb|��Xߵ��ɼJ*���n7J��3���QI����ڱ���ޜ������?��W����^�yt�=���ª����ǲ�����<�M}!A���#Ul�+��^Ge3��{1�� ��0�g��_�8�0X��?��Զ�bm���	!J�9h]=�����k��&?��O�d, ���1� ���6��a6L���?�o=U��2nl2�pP��h�x2��Gb$|��/��D�y�I�!#"1,��7H���9�T��H�A�j �;ί�6��v�>M�������j����c�$����g��4����-��x/H��O����"Dʥ�t@��q0D��5��?}������c~����#_�)QG���9q�}�9��·���ќ��z��p�!F��j���i+�z8������S-�	t�{K�a�3�YG����x@��n�+�#���A��X �?C7�pZ��S$	pySC�|%�+�� ^��?��Z�8\?LAG�~�a�!���k��������y��x��+߀O(��s2�����u��o\h��0@�2b�ۙ\������x��9dq �"ұ�x<��5+�NV��	�v�9lNSX�� �@7ކ�S�>��4!���7; �Q��dV�F���y��c5��d�<
�o)�c�!5}ݡ��,��8ׄ�_J�$�5�y����\��)O0Q��↤b�~K�����N^pm���VT1B1��!�@�R�_��2B	�e}��T��1/����8Ǯ����r\��(+ �5((�I�4�n����i{R���Ձ�ޚ%� ���*���~t�	�t� �sdj@1�x�'#���R��c%�_���梻��̀v6��Dy\�����3mm��u�"y�m2��?)�f].y0�Q a�8�j���y��ZӠg�=<U�փ�jc$SS�=��A�ǁ���i<�i�W�2��] n��ټ�T�h'���mX.�(8���o,����3߾at���Sl� ���X/3Fݏ�V����«����Ҁ�H���[��>��3c�.�/���0y`���?�s�t5���X�.���500d�1���[7[��V[7,t�Ǚ$8��y�gs�hŕbƶ-tiw��sve,C�^���!��7�����PX���)��9TƕE[AS�X������~	��3��;U�%@*f7�?�\(�����^gCۚ�$ ����d_Q0�'��>Q�ɯ��dC�����kD��?�vz��g��\��Ji�+:�z��x%�T��_ +�&�@9��2۰��r�#��_K�8�P��7��.�0m�w���_��/���'�e�Y�d{�䍜$gDQ{]n��m�
�s-@,gvt�\el�B��X�c�N�ݥ<͏����]��G��������L ��|�����$b�Tݝ�c�3��6~�dK�&�u�������ף�(Y_���o5_���7L���]�Y�1\��^�Ȟ�	ѩ,��?G:'��>��Ͻ?�d��M��(>o�F����YM���@"�'��T��]�e�Xμ<���R�� .m����X43.��im�!/�WGǙ9jr�|*O�|&�������O�(#��BP�����vp&"W
�6Z�#R�#��,v�-�'9K�q+3�C�wz��!�'�������o.���s��c~�:R�:-�3����Gz����4M��'53�m�&gJ��Cc?P !s�LL��M�4�Jsy�">����^��:�=��pѵl�)�:7?��,3�����b O��d�:��*�A	(�6�?xB"񤦟��=)^+��U��,�O��L�]<���D,����l�R�]�.7�����e��*Rp�<I�d`�s�d�I�8���|	s�xTz�Z~ .���I �:�e��C��%���	���N@�&��S� 边��N�r�@��n̡���*�F~�1X�9~X�� ��]�W���L���9��?nw:�����$m�q,��݋�r������,<��8�`���ш�z-���oy?Hm�\�<8�G�����ځ����3�+�{=�� N����n�N�� ��^5W#���5,�N4��| '�f� 
����3J�N�����E��.��%�⧰�q�E�߫��-���S�$bo�����G)�١),���Ӂ�M�bz�fe��?_+C�~ѐG^1FR��Y>w;rv1(�B`ڢ��j�ߙ݊6�e�g�{��~{�zTWQ�����*�G������kn�vLicU�?��	���r�zq�~a��4�8��CsX�w:��hR�z�8��u��*%����cg�a�Ȼˈ�D���b:`E�ϓ���*���<k):�g�cA�8I��n<\w��֤V<��Z?r��v�oy2�~wo2�W*�<�ꛩߘ>+��{z|�R �[��;��m��,�c�x��A�7�g�|�)�a�5b��6�p_��;������kPlOT��ln�I�nU<n����������`��ڊ>�ەG�i/�x뤒�/{��b�	�
4�q����
wE
��I�tȦw懟��Г[[0�nk�+^� �=bc��jP�g��wѬ�	���]�H����*6�C�>|;�����������c,��l��f�Оj�)���B5|>�����V������X	�)Po��5�Tb:؋G4~;A�������dc���0r�?��*t�"�ZÛ��c@�Br�vߛJ��{
 K�O��u.2����#ι�7tΘ5�A���$�?�������)�Iy�P#EAv�	����u�;"� ��}'��,*���z��<7�����T�Y��K6K��e�PE�� @��WbZ����� ����
ģv��پfXϰ�v�������ez�j`�B�~Em��{@4�Gc���)�I�u��ZP݇T۬2;vPOy���n�@pUzw@	��̼&��h����Dރ�wv��^�=)�*�w���� W{���h^-���Z'-E�|>�.CZ���瞧�/��她3�<�ł7Jk���5g ��,o�za������`��ʛ:�4������ b�q��/,���@��یi�@�k�$�: ��l��R��~P@�x�Ik�/{�ˡWd=��P�s�5����оy�߾�Kʱ*���}D�e�x�"���e�nO\�{<}m�zOm53q�MQ�i��.~��݄
�-�~�=����1:(���U1-��7J��8� �C�qO�� �0��oJk1(�g�(*߹��˾W��N����!.��a$�c��I�*�n5�BV��3#p���4���"&DT�@�c����q��66Z��>����P4�=��p���@�SF+ƨ��M�L�1��_�ts0�7ԐSEn�B8��?�A@"�wLm�V�ؔ.!��#`��:̝��������}���_��ڃ����.̑ˋ���ĤO�O�r��S��i{��x$Y������>o��ҽ��l���m��uL2�z8.Uc�D�<.L�9�caVg�( OA+�/~���F>�^{c1���3>���Ը��P`��ǫ	]�j6�Ԝ�w��5���ݫss��z0��8M��LT�K�ۿi�߱�r��# :���Ƅ�v���>5�J�R_!��6h�0���h���X��|$��b*	�M��f�/3���6���U<n�F��R���u,I4$t��n�
7Lyԙ�3�"m󤷮H���,��R��@m1�o/U^�,|j>��"8*�
M��hsaǤ�d���pۂ#��/��X�v�9/	v�V�kߣ۽8�h&YC������=��w�M�X������O)�[W�k�����,��s�N�Zw��!B��
/���v�J�e��ƈ�!��%�b�fmJ�j��xE
����7�M�J#�
y�8�c�\:��(�����T8��lM�8
 ���qv���@<�S���8 ��7��7�[�f(d5p������ϧ��o���a>��OAPcZ���`+�P�f/����? .w�ߘu��}�佖�祡h/��g�?}~���q���!�X\���iv�����M{���� �d���k{�����
���
��kl�Р�x ^�WK�#��0�`Q�RM[�@00��0+�$����<:D�d��vlˑ��� �T��@^y��@����i����@^�����Pn�3�.[pS� � س���W�hۏ4T�n�������gp�A:3���(�������d�{����S���ỹ� F�%;��-7w8y^(�yV�����h	� �ΑK����a<��Ǹ� i��&Ĩ�����kl��d��8���_.8P�jY�9�Ϳ���?	hh�����-pa^$@��x PD�aU�]��;�N[��]%���
�tpF̽�y=Bv��A�Ї��w�����v�;��B��u������V<�GZ^='�Y�B���D���6� ��fS��d�1��4���M4��]���g.��9������HE!(b�L ���ߴ#3R$Q��;[���_݋�E ���ƤV%y�k?0�� I[��l����3*b�pkҞ��h2p]N<��ɿ��Y�ҽ��r��j�p/�k�"��"ܲApĀ/ۨ�kSJ9���o�����)[:Y|7�P��B�6   ����?߶�򛰵���E�J%��qb��~B�/Q� #p�4qo��jİ�8�F�1XwOe���z8��w�̳��h^�^�S6y��C�2�
���&+P�Ȟ��K]�.�U�fT��"����0MlCޫS9aX%0df����`���6%�:X�B�lO]�ƅ9uo�">%��T�ȼK������Fm&���S��7��E5�/3��[��:��c�/�`���/��w��L)r.:%�V|�n�����z���������mt�^���L`�	*il�
q�n��Y��nĐ��xc3��J���n��b5
H��'ɛ �Oype���%�,Q�J�X��R������5��6�TÃX2��?�����R	�d3H/�^�S6*1�K|�}h�vԭ�R��c�7~�9���Ak\�n���>{���m�Y¾u��.mB����]LyL˨w\��?�[w��/����v/���`��"�d�ҥ�P�����e����q�?��0̠?�[��E�1�p��@��]��K�w���.t�f�&IoK����g"�+[V��5�����<t�y4�d�3�b�����uK[7~���k��g�2�����:������w�5� ��G����������������_c^3� ��J�y������_��E�ڛ���6��C��%�O|<�oז��r���,�?�aO���6֤�˒]�s�C���4�(�ZG/&���X�:�f���-
3-�R�I�W71���v5j7��਑Þ���C'.�B^m7yl��{�˵?�n���,�����9�ܽ[�s(�ȏ�<�Kcm�I���xfs�~����~Y��;���c����.�E[���(��6���y�3Pcs�#rq���d�0u^�B�����}�����7�T��p���W9��>�P�W#�R��af�o�,� vDxs�waQwi��o�ǎ�m^Ӿ4<�D�{�9�U�N�ouj�sɲ�VR9���ț�6����(K+�e8e��k�7��n�3��BԯJ�����87�x��D@�޳=AAqHG="��ȏ����uQ����D��d"}�^�cs��n��)�:� �%ϴ�:�T�4=�4t5�ƶ��|���|�g��w�nZ4H�s�^�2!��O�<ʑ0�ԭ8��-��iz���mw����^#�;�x��,/}��qm3�����j�!�_jD�߅Eg�SS��jc���jsH�ѹ�Q�X4��b[0��#�?D�&�of��KM]��G1;~���s�~Y�a���
�^>q��;��84v���z6��3��=���59=M�72���h=��j�9B��&~wM��U�K	���ٵ*�g�W��v����V����̬Y|��7�.�vQ�'˄���G֙EJ���?�L͐]��^@�+���;<7��a���E�2��w~"�c%����ˌV׺\P�((��'�r�Z��b�l�߇q���qo�oq%�#��=S��2��v3�J�A�!��*��"��q�k�ʬ��~#���<q6�@ڙ� w�ԁۖ�{h0{Ű���(Y���oRE���;[zyG�z�7�v�d������p�-�:m�҉иk�?U}׌�D@n4!���Tz]+
��H���M�d��u��J�E���p��i�_Z7�9(�9�S���l@���Y�ny&3,�-aZ9����[��p?�y�,v���g��(E�%�?��k�+������|W+!�|x �5�N��'����ŕb��Q��B�.U�]�2�������7�!6D���9W����lH��j��Z9�F*z�85#ńH�(��4��?��ѽV�zJ�k�
۷��*|KU:-�D��B��|��u�m�󙀳 u�,9�9Z0��U��M���R��%�&4� �	ŝ�|�<��*���:�ۼܑIs��p
r(�ĸ�몜�mb�W~f��>�/e���A55�$��¥v�x?Af^�j�Q:lKD�XR���V<ݿ��BP��tQf��a�J�����m���
5�ʖ6��I��BJ�Ⱦ���R�P	�P)ʞ}�[��k�dwqm�~���]���<O��<�{��|���y����o�6�6ba�.9���&����e���0�Z$��3��je;k6�Kl��X�?����55�ܥ�«'��Kf�r,W��N�i���ͷ&��k���L\�����7���ǲP��?y���4�0�D;���y�+�#�����ƫD�:�X����������Y4F�Q�J(��;�j�����M��-��:y��qb�a�H{߿�o$�+�KzM�-QtM��w��n�Ƥ�5��UD}ll�b.�Ո����kRZ��P,�2��L�sơM��U,��D{�� s-�h�;��Y�c�H�"���bQ��;�,��j7�5ʻ�]�w;�/k��wTM�L�s��zl
��t������] �K�S}��_T|��ܓؗ�1�dd���?�=��Mm��ء�T��5�(	�Y�@�i �;S�_ؚ�!CT���Ua��&���°��:���S�h�Yev��J�Vx_Ul��S�!�Ff�vOms���4�ԧ�Ш�9�a��xZ�X�H�s���f����1S�cv��&ʁ���	Ղ�>�Eɬ$b��U1��&w�R|���n�$ߪ����`߄�C�� l��&��V0p��2-f�|A�W3������+Y���J���Ҋ�.5��=<aLq:�v�Z�&u�~`n>�i���Ǆ�NF���XV@}�����j��)R��U�ַ�Z(�r�}�@Ǽ(_�x����)�\�}�6
K�/�:M��p���L[�H�C ��oQ�`N�V��\�᳀/AL���wiX�\��V�W����"L�S@KF[�\ �%"����/xQ�^�$ `~�����L��<M-�HqMUZa�������V��\�k����u}=DQ����~
B���i�A�9�����b��c^�	C��l�VӍ�t��rW�8�~�2���]��d�>k8���]�6#��YHu��t����^���:9c�F�^ڤ _�����hN�Q�uu�h�����¡�R;\�2mc3�F߆���4�yg��H������s��<�,P�����W��*G8�Ԅo�ų���"O*��e����eq��KDԈb~8w�kF1{��;/�X|q�әj
?�����`m�@@0���3�7��3�	�b�����_��������?3x�1����ѻQ@Z�(H&�Kз��M�n��1�����|�L�˃E�8������!'z5ج#~H�w���M)�u7�7C����[�'o�����uFSs_�`jX�d"
��P)񒶷��///@d�Vb
��	ӌV��`�xn\�^�C�<n���t�8�4�N��Y�:�W�Au��ڝ�]�R��)�jX��sFU5ܔ�W��Z@�IĹ�Cq�\o�����qV\�܆z(�9ځZ9��*�c�.G[����`��'��F59�A�Bt�����k����fYi�޹��o ��U~4#-�N䣘�R�͊Z�,�8�HG�P���B�,~�V�*A-�S��و�4Gr��o+�~��v>���%p:���[����~I�VB��y���Ft�F��A�L����#���l������zR&i��+�O�����@\6Х�xO�ʠ�"����pK�6/�0S�r�罺§w2Z��k�n��!N�u�x�W��(�W&�������6��P�t��f��<�����L�����z�<�8�JX�\�[��;���쮓t�s�U�4}L���o�pܿ1��Y���[�FF~�x��4�6.�l�������x����Jt�v�T�p'R�@\��g�@�x��f���z�F��y��A�1���;�j�%c���v~�����{�~�M�YOR��S��Z�	#\�"����rfh�}�hj�i`��oR��6�Eʸ�"1�ҹ[s96���$��OZ~Xx���I+�p��;��V��g �`WT+E�b����^���Fr&VH�*���|$��b�I�~JPw�#e��Rh�\OT\܁��B�11�j|��1s�rWtտ����>@��Hpz9�i���U>��e��dĽ 	NT�fƛN0a�ʵ�j���c�fO_(з:�$F0n�*o!:5!�g�t�%_�[�ZLe�ۥ�c�rϟA}���-�5��/�)��1ȟ�rkc��V?v
��+%�G���H���&��(d� H�F-���[ǜZ+��YX"T ��₳ ���D����!4��K~�LA�3lf��$&n�gd��k��,V`B�������LOv�1�uL/1q~g�V��yP֣�������G�� N�X�Q�c��@K1��+�A�-O�U8Pر����y0`:)~��d��N�>��fe��k���FQ#VyȂ��T�VP��ll]�!���u���#��x�Z�fy�)D����eȮ�a?6Y�r�.4���C�iὂX�R���?���("?�~���S�.G$��o��y���f�5����:3SZ'ԩ��פ�b��6h[�ܶ��3�f��At6��(u�k�� rg�.i��E�t%�ƍ꜑�T.��>�H��s`�)�En��tN��Fu�=4'��8��*��4���\�>��'�y,����F�����Te�y$G$6�=��H!̈́� �˜�൘����e/4���jZ.��˅p�����+T��bўˡPM���N���yw�����
Uq�q�wW��C����ܿ����#�Ν��@���h�񕩪\�D��
��eo\ܙ��Ƣ��

�6�b[Or������I9�6�@�@�����@�"�7Q�y6AVAf�ys�㞹.i>�;`�(�q�ڍRMd\ʀܨ�2�VV�Ke�����SK��{�S�����d		�ƙsx�鴇��-�ɼw
�*z]�}����Ź�a
��kp[��?�Pe2r���Y�
��f/�!�z1��S��PX�Aisb7����?j�z�Ĺ�@�,cCn��׹�������`���Mqǟ|"����f�����2�g��^�s�������b��/��M���8C�- �̯���Seݮ�?���?B�}�_��{��8���  �����6Y��ŭ�Q�5����\� lg��t^��L��$�)�|��:�fj@wVBWd`�g��U�hn��(�R���� .gR%��Q�O��d�~�����`?�ȥ��b��%�tDN�\�dOߞ����ƙ��ȓ�����������:����"%�ڢn��I�'�F�.w䴆_������\�����7�G�#C~��fr�J�:��u�m��{?<e��jG���~�vm[�zltA�X:��j�s�nW�Fr���mɴ#}�ewI�k>�a�ϻ�ϿGn������Ѓ�;��K�^c�I1�G��h
,%�k��\������( �le��\S��ڭ�'X�����&�2��%�FY�br7�|�;���L��v�p�&��#�'��Lk�O�Py����;z4bXd[��̞�����+9w���TJ��'�1���Rp9�:�6��[rw�?��G~�W�W��?Ż!FԀ��R�L�\��Izy*�ea`�)�t�kBN�^69�a��Q�n5m��skc�45�R�n8�ޣ�?�B�3�G	���$:Ɲ��e�Vm��'g�<'�^�>���ѷ���9E]ޢ"�[��ߠ|]	�-sɥ9��$�ǫ��4��3m�R�'F�'�:կ�4dw�|���[���P�)�T�CJ�]���#��[�k�C���9�����	Gth���:�s�Ĳ�����XWԃ<V{����ϣeiN�af�w�\D��������yH�� V钰>�C\��� �Y(�Ny�@�9�XE��3�x m@z���&�"��]�Y0�p�c89�\���Ε�O|�*^�Oy��x�a�l�	���i�S�{A� ��������3o�)#d}�\�r��#�Ȭm�W�vPf3�A�	��0\�G�������Ƈˡ����Y��S��n�_��[�d�jy`u�s��3SN4�y�Z`��R]a����|���xJD�{R�/���1/�*`�1�����lk���5�yxo%�tU�� �S������3��FHص���h� c'y��������ӌ=MPl�;i�5V8)�#|�"�떳���{h��;�v��bg���� t��,�K�B���ˌK�Z�R���܇%��Ʌ�:��M�U��&�!�"���ܐ���U���_.�--T���ڙ��,�������/|A�kתr���l���>�����̛�S|���©"&�(�:�xK��D��iHH���R��n��a�=]�����_>��j�����>,����U��|�{���x���O����t�:ک�\����	{���� ��>c-E�qc��}�������KߊƇ������IqI��V��V�s�2���߸�s��Fw���jIMߏ�s�Cj��������*�[K�[Ϗ\��+We����~�ii?�,^�s�БQ*����`y��i��|���k�v�C�iw��3�o����:7�Td��q���5��}L�.A%���<��\��������:�˻17�=��A�(���"APuߠ�����4@N��UQذf��f��S]6�y_S�a���"9J]��Sk��*\�Ȧ�WO3�awid�hR)���L����t���Ɖљ��<���������B�!19�L���ʬA'/�cx�{���j^{{�!a����
볖�)#����W�Nc_�R�W���a�A:b�̐oκ�k���A���[ŘR�`��s��l�֢��"�q��Xg,� "�-�,�&�e�2P̡�o���8�9K�e-������ľ>� dЌ��]z�5��ؐ��!�7��\ʫ
�0q�[^|ѻ@$��}+�ڧI�;'�A'�O)F<����_�~�T4_)E��M��>~���0l�L_��pu��9C~�����Gy���\����ƭ{X+ٔX�@���K��,��Wb;a9W�NhK����*���'�;b�2&��_R�.'ks2r�56�˫�;�5#��G~w�֡6�B2������x�
�ƒW�=�b7�ڽ�J[�5H���&���(5����>?�4Vh����{rO��d5I-K[��ܟֲM�7������YS�A�Aw�+
o�֚j�na���{|��}�6�0���&��d�d��q���CaQ�~��Q	Uf��4D���{vŠ o�1�'
i&�.cQ��n��t�o�ʉ�O���(���ɫ�63�4*/����~�f��%bS�J�Hj��{4��v�Q������T��C�Z����Vz��0��-��P{�֥�%����y�*���j����ZOk��~����jk�А�ֈj�(@���xv���H�"�ܙ �=��)"_1�,���q�ڼ[�|kA�\c��]�˃��_����;*�z06zȓ��<����WŶ� �Q��3q��$�r�M'Yo�VQk7�zSsF������\�'̗`����_M:RY������n|s��W1Nt]��4�K �)�i�*������'V�#x�b:P��������	M���P-;|�|�j���lF#�>��}�N��iY��%+�/bpsG���w��i���d^�v���Y��	Z*Nr��~<��D�^5|�e���P��'XN�[w�{�>g���jp�*�DG&*�N��!�����z��	T\vm����c׭ڼ��|�� �zR��0��I�`6�y·1�����3���Ip��7��`
���q����~���r�����X5�g��9k�ņ���o>]�Ҫ1�3��gY�n�"�19��6��F��*'�_�>oR��%�K?�yY\Ԭ̝i8Ծ�OcP���}�W��m#������|����T�����Y�R����wc|j���zF%�J��;NNUe	<��L_�$l-�a�iy.T�H��Խ�N��]z(!y,]�1�WeP��pV��>ڕT�١�HG�hܦ]
�nƒ`�	t�\/�,�)��l��W����%E�c)�E��h\S�k�a���̛��Z��Z�xd3�P�mq���Nr��Nc�A�c˱�,�VJW���9w��@ޤJ+�]j�Y~�R�㢟��C��9(�!I�_<å��p��3+ߣ�!���q�H*Z��jM	�h0g�%"*�(͉�$R�s�V��{#^��^N��G�r��~�\��3b?ΨKw���HmH~u��U���5�5�O.r�]������,E⨜��g�,�%�!�ʺ'�+�pn�×h�D�w,PںI��<���H|c�%[3J�|;�����\gnR	vJ����V�H
�6#þ��GoU����"\'���S��z"���q�<܋��T8���`�EzHQn6�:&��C�͖lǆ��O��ݪ�����y�l���W�-�޲�دrq����?Bf�0���S?��P��9�tD�8�}��%���q�s9j�dɃ�[�X�������P݄��.�D��EYM;��3��ѽ8���#�����Y�PJT{�x3�+v7JJ�����;��5���g�4����a~���%=@朗,u�w����1�MWŮ���ѕj	��
ot�>
eDޠ��>���-�����\i�}X�hWoIR����4�H��L㋏�Pa��3�r���7y�0�G������2���#%�����*�3��ɪ,�n�H>��[���1���El���������R��Xy��":n���oo�wN�\����[�?E�xO�ڛ�-�פ�W�D�MԟmQy�3pf�>/�l�A�x�g(�cz6}�2��t�CQ�� ��VE/��D$��dGN.��z3b��Y֒V�Y/�?�����Q�t'���Q2�\�
戤/�x�'�E����;��q��G���1.���9C�Zu܃,�W#��䯏wU�w�����mZ�
�be���O�i��{�&k�\�9hK��y�S�X�&����8)�<!�/h��x:���#V���nbuZd��|
N�E�8�u�N��ب@�xs��G5�Q��{/�b���r+"��;����8`�\�M���'����4E��hSo��o��{9>�-@�x�P̳��1�S�^2i��,'�[0e9O��cյ��ɾ�T�݁��(�-�����4p����5¬�nH�䙗F�e\�Ëw��Ji��������3�u�&[z.�VX|�m�;2�pN��&bH=�)�}�^������5Jj��2S�ac^��Ɩ>���?	g��C3�A{�5�)=�F�5Cب&��V������D�L9��k��4��=<Y��Ҵ�)G��)u x��ވ��>��.C�L��!�4b��7�Du+-� �������(�<^�h���wu��?e�v:��|����v��>S܅~�O�7����/ѕ|ƺ�;���L,w�z�M���D{��]Z�i.�J͡�������x�}E�Bk4;G��ڏ�ʁ_@��'�4sRyNM�u/�2hAـ�[���e�Zλ���}l�e0W�nc�WY�@ [�9)7\ɜ���ʊ��K�ca0C�E3$8)g�Kb�K�$�h=]n�=(�<�1~$�u���}5����u�ʽ�BAW�t�8[*�k��I�ً�Y�����R��rƸqo�s��ƌ�.l��KP��KާB�����^UCN�E�)�rhE�u~������TM;�`Ne$��>*2 ��k.E�E�8Xd>�7��ZaS_�M�ٿw"�B)M���k?HL�yW ��*�5��D�L�|l&���N"Pj.M5���2�X;���y��M��Y���Hޑ���c���j!�Ŋ6	�2;Fms����RA���<$�/>���r��ċ��H�r��dXT#���+2�9&�+~�c�0RJu+(sX������a���J������O^��n�W9�l���ف��w�_�tA��Tn��_�m�x������#���>��[���y�i�v�Gh�+u[�>V"r���4(���q5IMVYs�%b��`Y��r�;vX>���V��dx��`K<��k쟟S�s�Wþ�3� �Hf@O��Vw��U�-:����)�=���c@?��Ar����n���f�pN���]	��M�cfr'ܮ_3�5-�U;�;��G�2n�Ug^��䶴�/	KX6D4��_p2�s�C���H�J1�����y+��I��~�H�ے_Uu��*D }柿	�C�w�� c�̜A϶b:4("a�{haU��B�C��ϵە�h��:+���;��@FB�����G���]�a�(�����vҼ׊F������?�Y����ӥ;��ɍtNZIN	���#S�C�V)�B�O|6֏���E��U}�'�rx��ǞO�Q�;��u`]�zvu�E�p-��������;V�׊nbM}@S9j�,#��V��Y��:vGMџK#}3��b쐨D��b�u� �ʣ�!�l��w(v
^��QH�����=yKV�� \�I���Q�� 	,��I�7SX�Kg��n��Qуd�����R.=�V&�u�:	9}+����!_6\Q�cݘ�O�Z�����b#��b}�\n��t��L�帋>5�ƴ��p!�5��*��䰺#�T��`�2�<�b����1�s�-|v2�6ND?g
/6��"�h+O���e��˒��ZQ���-3?�9j�ʑa����1���G[�`�m%M����X��=�s�nNy�����v[��z[��*��T�����lE�T~��;�KP��%r~}��%t
 䃆��!n`���Vڤ��r�י���; ����ٲ����-N�F�\s�I� !D���;�'�0���W��$�6�vG���
��I��P������+�o&����N~؉Uў�?
'�,&��V
!xՔ�'\�dU���X���XƱ��� d�6֠�X*�E;1�R�[R��ȹ�g��f�![���]�D�����εl¿�1�x�X|NQ���꟧��-M�!>L�?�|?2\��G���L��k�f����;~ћ�K�I������^e-$nWv��m�鶵q_�P�����'e�<�I�.;eǎ�-{C�܋H-����e[�-�Y?�	��v��su�����ׯ����Mc//�䱗32�D�>]��á1�h����H����G�b��5X�3,Y�=X�/����Q�Kf�0ӭ��e����W"��z�ܟ���Ũ�I��p�����1�t&j)��^��E�(^����ެ=w�G�=�i*��R��-��E��}���G)-G��l�B���<6�x�����~U8��C�pv����S�K����`������--1�.�K��1�gPfa�V�����53= 7H����)vO�sd��I]l�k���k5�s�%�w�t9�B���Y�[��l1����ɞk��ac��^n�A����7h�blV�/���b�V�?��>2\8�]��Q	Z�s�Myj�ި���b�D�5�Ǘ�����n1����$9/�q-��w^z���Arx�����ݳ��Z��	Q���R�q�z�"Ӹ���h�HwU�E�?=Ό�;{����K��:Wáq��F�L~ɒڥJm#�����s��|����࿨r�ԝ�e���
1��z�uQ��{n
m��,{�fyF�d�r���1�0?�����]��EX0O]��{K�x�ci_)�⺱���k�,f7d$Jԭ�����g�J�D��&K��nرn��8G�Q�M�u�>�2� ��S�e��ײ��X��]�:�?,F���N�/H�xL,i�١��i��ҽ��L�53��]�бīt��T֐�����̏~U�Ut�������=��}�{g�p"M�t1�D1��W]_�?Q��O�/�R���L�nmٕt�p�*�Rf�JT,���� !��e�0����e����cӺ^m�3+���?me�*��+N���? �e�1S]#c���ެ]���d�K���Xb�Y�^�oWr�x��쾞zeކ�����`��R�j�����e��J��i"�T�v+���%�-K��OmȬ���q��䑒�-J�����ǘ#y��ړ�9(���a�Up��.G�L�.��h7X<C&���11z�މ�߇e��?\�^|�l�Ē�,�%.���G�\�X>�l���1�ǃ�ڄ�>C�G�6�z|��hG��<���_��U���e���B��dk�B)���YY;����VpEO�:ñk+�[����FO��'D�<�wk�"��]�ٟ�1@L߇n�̜��qv�p�55�@�Gߓ�	aPKC]̊�3l�Y~�o�3^o��T�ڔ~I�T~lm��T����xM]Y�d3��w���n��.l���/���8vo�o��)�~q���"
O�6�=�h��|������Q��ީ-�i��p���zv������F���npa�Д��%����w�����-G8��BT�1rz)�@6^����՜T, h�u�*R.��ͯ����A�i�n� ���.}���6��;�dY��4d%Ir��7����t�/�]f�����z���-��?�|��z�2y.��wh�]ea�"]䬭�����$�I���c��ĳ��ʭ���u�7U����1f��W�V�x�DA�Vo�,ߝf����O��7c�뼄��o<�=O�;�\��K�>I���A#!a9��SC֮��ȇ�����tؼ��EP��
��nj�+;R����H^ogo|�4�A��x�ɬ��R�&_Z�쫳��������H�}a�ʚR��"�t�ȇ~ZG]E�ԟ	K�����s�ȑ��"�Y*�[\�UHF�"X���j���A�R�,X��3�q���*ƒ�p���U*E�y^�$੩�A;�s�;Ѯ~h�y7j��� S3!6s�
��M}�c��Qʺ/݌|p"���fT+����9<&@��*�Ƣi�l��`�w7Z�(�C�{Gl^����H�%��c�>{�׎)'��!Ə��N:%�s�;W��63}|f 8y$�F��X�%i��m�j�xo��+MG]N;N�eo���Q�����!x������ʦoK��ܡ =%��a���;:��ۿut�������'��q{��;����*(�:t�W俘��q>�??g��h�=?�&c�P�$�w�,�Y�S�Te�zr�*ƥEa�8��}*���u`�m�I=�g�n=�1��p�OW������k3���O�#f`.R��h���n��紼�L��>M��|Zs�nތ�%�����57��c4�R^ 3��9
���37��oEmL�!�^�(�tQ���!�E�#
$���]w���N��V/z���,~-��j�� ���ͣ� g�͔̈qD�nQ����á�Mj���j@�.{�EL@mм!�1EY�MS&"G5�����85���tՋ�¨I�	
�پ/�o����9YǴ�r��5�{U��>�H����1v�-('���o�aKs�`��`�E��r���m���t���[��ln��)��nW�#c�Ò�Egѵp{�ô��ؒ�-��zܢ��'@O+�Ǐ�����TmEAe���n�L����w�>��s�����G�\!t������>�!��ѓAU"���[f�*�Kq4���1M���,J(o#���E���eǦ�)�8O+g�G�OSs��Oj�,iG��x��ސ���૟֓de�OY��>dc�2�bÕn�U�tȊ�Y?����8!��>M2�_����K^�{����I����Ȥ�FW9Էױ!C4ҷ�,u84��u)���}�[
6a���{��vq�����)əmb��}��r�ec�HQÖ����&�ǅ�|�4X�:]�"��p����i�<��U���lA4��p�Jb���2IE�
wT}�N�(NcmgP�Y���o�(0��0�Ø�|岥�=�=�|��=2�xf���{:�����C݉�g��RM����yG㝨ޅ��ɼ,�~8��	����9A���"��ݼ�@L�!���˝�}�}̑���hɼ�	�`g/Q�+�0�N�<��Q��m���{�|4j�
���l<ґ�!�yd�>�_xR�۞����,�,Ag������&HB6��V����IGbo��gz�l��� UXp�V 丹��cp`4�E�͋�
>����`��5���6���<��>@�@�L��
��[/$�l�Ó$�5l����䵠�[�,�3� 뙷n񖎋����C^�4u5ZR6*�����?�B�@ �.���_����H����N��w羨�bb����K���O.^8�����p#F�]�J���""�P��꬗�Q��Bv|��1(j�R�dM����!�\����&��|�H1I��X�ՆЙQ���K�
m�L��`��Q��V*��0���K0��Dex�XCM4E��r���J2��n�{��K����1[Ϳ��哆��M���b،f#�6"9��.�Ab3�K[b�d>�?uG�=6��:����Э��v�U����NI˶� O�ݱr>�O�f8y[�ЀL���c��T5�g�W�Xo���[p'� ���&��r|8e��,�߱�� J���Z�j\Q<@d�8����ӷ��"�߰����h��j���Jl��˘��}V��S��8�`vRu�L"f��_� %d�%Ǘ�+�[��r�����?;:��4GE�:'��_����O3��ġ�	�\`��[a�ۖ�R��� ����u���&�0ҁadpI�WZ��VڣfM��d �䥰����I	��mx�1/�����G=�"jp��`� ���Qu��U�W��)f�����а��ݻ��5W�A����ڪ(��C��+���4|b���TϞ@'��$�`X]
��--ݝhg�v�����VS�IW�Z�w���V�:�ڋ��}
b��	a�Ӿ��.\�I�q�t�`?l 7|�&n{��U~QF��*���&[�,r������=��]Wj ksw��`�y�a��3�9�b;Yf;� ���O�	���1��W{F) �g2m�� Lm`m(�ci�=z����Uzz��<��?��䄚�Q�s�B��,���n馘�{./��[l���u�є���d/�KN+�46��jW�*6�rM�^���x�5z�bG|{�����`ׇ9aǜ�G]��Ū�Y}�.��6#�VSo�� �#��M��r�I;}A=�Q��0v����I([�����A�k�hVD���]��1{k���M�:}����lR�y���AA�u��=�H�����,(b�̺ӊ�r͞6G�(����A]�o7�n�b̺�e_�5�7�I���;��#��!�-Q�ަ������(�{�6C~��m���XdS�\*�	ˏ�(L���_Rs�\@}��`X7e�/��Z�p�yшF	T�HП�d0!Wk��q��P���! ��M�����	Eb�57E�����f�[X1j������&�PY�{ڰT��Su�䞇N�c0��6��>��l�f���L��a��@����N�#{�v��[!8���*�;�DΕ4�hU�E|�C�T2ѻ4V7�=��°�Ǝ�)S�d��G�GЄ�Xs
\mƭz�%I���g7�~9�܉O���-	`>����h�	��:+1Ú�@R��I Q~��?�~Is��e���;�ݥU\��9��F�A���E^�.�W�$�[�¿��2r~�J�;�?�:!��	A������&G�Qx�EIZ.)���`/&خa��YE�r���&���eW�7 .�� p�� �@�t2�n�fy��+e�«;
u7��$aW��p���BMzo�K]����g��T"�P(v~�z0Mw'��l��o�!�X�;~"\;�N=)�+)�#�s���2��<�*!����Y��f����T�!04�{J�`,i�����B'��uL�@���~f�L!��&Ͷ{x]����-Zs`���l+�
9X^��5�\��$���?�Qo/
�] �q%WuM����~eG�^�f��U�T��qƑ2%w�ى�J��tw.�ůK�]�#E�-�c3/�E���9U��̫�L������|��"P���B����ECڜ�#�N**�l�T{M�D �"�U��j��m�$::���~�NA��ċƨ��g_^�|�\��Rۿ��9��#�2Z	!��^M/Q�Q#��dz��n��f��� �%�)Pv�F�Xj��d�O�b;c+��0�ՠ��ler�ho��*����#S/`����C<KG��Xg�`�#��ЮW^Z~��=��6Z��{���Ŷ��2W`ji�ԵLWյ���(.��ۘ���h�`^�׎�~��7߉��\�"&Ѕ��׀���x5���WM�ךLAޡO�[�[E�/[�cjV�.Bf�6Zp5-T�̔�""���w��8�Z�E��a|�*t���v%�|�v��I��z�
�،�'�*�EO#�<��78���{�Vr��7t@�F�\`�Z�_TE0@�i��w��/�
��B���2&|a��ŧ����W(�NY6;µ�R�a�8��('�#a��ՂH���� rd�$�2�m`�E!��r�%�6�})�|_��;�
��'�[�#�!d�~��R��\C8ƺ*�~��`߹~��6��W�
r��&�;�Ծ�\w����/�g|����K�ĳ���~��t�ɉV���/��=����@q����v�������i3�w[�o��-M����5-h_����3:���p̴����i��ϥv�XT'� �h?��x���W���p�k7Z�I��4lc!�X��x3%�-��Q�Հ`�F���������@��_����l��By�]i�a�=iF���,�h[�*�D|#,��y����̍?���dV�ykߍ�	6��b8���A�?7Zl��$C�������>8]�g`��}4~�}V�R�K@{�k�TT�?77Є �6�fʲl�.�@mxSr�Q�xIL�Ƅ��M'�/}�r����X��r��iR'C�6R�sP;�aÇ�>� �0�{��P;� X���&8�E �F�n2�蒱��:L��@��u��Ƭ�:��������v�?������F�`�N��)�f�<N�)[5(��ϟQ�~	�"�f�(�V�-�!�۲�c�+Ńl�M
n��➻�taq�P	Ƿ�@C%�moڠ�t��U
R޵�.��{�t��&V��;�G=���n��Kͣ,i�k�YIM�'s���R�{A�V�k�H�T��~r���&T��"���%0̴ ϥ�zݫ���x&b�碦v��~�Y$Q}4�v@�q��ǃ�-o�����<�P]��ź�`'k]���A�!��D+�]x[������;<����OM�'�3c��ı����Cs��h����ǟܹ7XȓrX2	��,���%� .*�q8����� :uO����0R,�;�����LN�6�OpĶ����>��2��˝�tKf�:Bg��{��J�T?͉�Q������S������0���C4�
�Cc�7�y	��#�{Ba����/��x��+���k�Fy/i�`����y�DE�A�1+�mBG�������+�|��H�R��-w��.�u��?���B�YD�/�S��ʜ��L�{^����3T�?�/�.GI4wd���ೲ2HB���4�/�ލ�����%Y��Gɀ��2x��7T�Zi�s�p(�A*M��0
�n1<5"�㴥q�� ��)1��]>{��$ġ��5���o ��<d�?ZD�z�aDz�i=�6���?R���4�Z7�`R�z�z��:-"����}p�3
�������i%xe�E8�A��/6Σ�-�_�������ǟ!˟ݩ:�l��Ʒ�]�N�ѭ��\[UN-���
H�W���_��֟Ӱ��K�`��0n;��k	��oCT���X&��[=.�<��������$�zal둂-�^�
3�2�mē����O��a�v�T�ኘ���v�?^���o%`j{��Q;�r~!X����MҚ�!^��x_��A��m�?��~���-�p�3����N��)���C5�I����-����a2m���_J_�v�m��p_����K^����͟;���Rλ��T��ol�uc���S�ߔl/��V���'%�cMsCu5�.Q�3�W��$Q�8S������մ}��T����߆Ҍ����y9������=�7=�n�*>�lC��6�۸�6;��;���-��޷�bY6���Uߖ���H����0�'4��#�W4�R��r�f'�_6x�����t͍4���E�zd&�zتɼ�WB�G��}C���Ux{��K���9��V�#i	�3�
�=�YV����َ�$�{�3�-���
g�kG�o���Ic���	��&�8�g�����xF��R�2d�˦���XW>v�?S����TZb ʟ5��q?��m&x)Ӎ��9�Yκ�E��Mv��7�+�� GP�܎x����ʫ�cw�.�2��&�7��+�g�<�h'm�w�8Qb�S�ė�g��(��p4���zd�a����=O�f�C��L̙f:/$U6���������D��_��O�zw���
��H�9�>�'.��Ĩ�A]�y؍ʕ�|��ɒ�Z[��(|{������ξ�����#�ʡ~��[�g��K�ۚT�t;�eKY)f��yN�}�c�B�?��2��K0o~D�y���Ҏ��-�z&kx�"�2�o(�n�$��ܻy��=Lz��w�??Q�U�~�j��[�E������-���f]x)�}Ӗ����@������'"2�û�4�3�����XbO���[ҭ�\HԽ.Xm�}��07���T�~��k>\0�����?[ұ��<���*9f��L�ts6O��<W���~~�e5�M�L�0'�'��ue_�m±'���{�+�FZm��\]i $�6e��x��sgG��58���g>�� �^��w��>�
F�����b�0]��:�:�:�O��ι���Bp��֙���@e��f��Χj+ l��g��,�	�q��)<Q�#}Z4 b�K�2���nb�r�gs<[���������3Y'�-�*�pG3W���=�7���`C7wu���\X�YR��e��$��p器ù�&):�8�iQ�&������z1���k�	�ҕO��t?��� �[Q���m��������=���E���:z;jEe8����[/�G2��,D���7=��q�rp����l k���U��d(p<V�������ժb��X�C�\�i��B�KiGfs�C��@<^��bϒ��7|(bS�zq��UE��k��@�8�Ù1g��<� �ZyU_�V�V����P��b�zp�����h·���n[�M���)����$�qbh�r�y���DW�G�N��u��N:|����4TK3AP�dxV�GQ
v8C_9~���a�L+��N@%)�%<}��%�ֆ�5�yBz�wo�[y�IEa��4c0]����v{!��ldĸG�7"�lL��i�Е�����8�ȉ��6�m�� ��J8�>��')n�%�����r�c�:b��<�^�}�R�#]�ie�I��HGIԽ�� ��+��	w<�,|L#�[=��������K�S�L�S��qEd��7��ᛧ	���gx����1�Q`�u&�Vփ�I?GͿ�2�}��7:	�"A����h��BH���A_�<g�ee���>������;�(К	b���1�p���XKn[�F�S�{���_�?z���8V���H�zQB�;�� }hf��{x�t�鵛C�{:[;��@��Ղ�)=�G�#
e�'�{ծn�=�;�d����pt�'��>���l�8�4�p0Eܜ�b�c�����g�/����eY�g�����wW}�Y��]��;A���C� ��˧.�.wJt銔u�T��2��B`�����؟���k{�ڢ�ޥَ������eVb�w�����)�/�O�5��?�z�"�W������{	��=���?�x�1��(��TZJ�V7�v���M�O������K�i�rs�9�m�>	�̟�����&���S:	)�e�I
��iяmeO�Μ�><�'u��ڊ�=�Y������r�F� ^�*������>P[b��2�
�<F�'R*��C��s~t؊Z�&'������Vҥb~� ����9s�#x'�_����\�-��@\�W�k��9�D��j@G��VkĐЋ��~�Y��v�����6-��8o�����Ȟ8��	m�Ԗ��_�0"-O7/�}��6�g�"�4b/]�0>q.�RT��D��ƿa/J<�vQm��%�<�g B���������GB��ľ�ס�]q��������g��eM]�v���~:r��{Yw��4/I6�^�z�g~!�W��[�w��`��>����r�Y�z������>��p��1�'M��eyʊƶ�A2���R_����_	��P|�S��љ�C"��R�B��$�3���\��ů3�.N�=|�T+FAd�B�6Xj<c�����5����{g��D���@�K�mpeM�g��W�< _�+�JT�u����/���lbn�m����}���n����g�m�����w����)���i���"��B'�Nԫ����WY|P�'�i��'t���w�sp�bh*�,�2h&��n�$4��=�ljm��( "es����^�]ׇx٨9� �/: �q�#�?I��f9]���ȎK�%��",�A�d�5qH���/�E"�E3`�]�)k:k
��l<q�ϫ����.�,,M�{��6B��#�yl���>�M�>�*�HG��ͷ�͑v�d
�/4���ׅ}C©O)��R���/h��/��^P�Y����f�W��F`�$�z1�:b�ˤ�s�ٿ���VÒ�9��b��k���_;���ہ*�
���*\*q��uRz$ބ��:�6_�}W�f���f�g��:�g��I7��{	E�Űj�ֹ��g"2����!ߜ�Q����k����S���	{�菸�����~�|�<�u���r1Č������Q|�7?������Ū]���m��3bg����-���9�lBBa�������=�ePq&A�߆1@�FPG�[�G��&|9�J?�&(2�h;�/�����޵�hO�f(���������G�&i����A�>�OD�+QVd\+�q�T�L�%{fo��yCƥ2B�#��<�9���_�y�����~���sι[{�i�7l�R���m6V���Ϝ������ąH=磨����T�c8G�A�X��LcsS��Sr��1��{���Dt�A,��u]k�ZW���;a�ᔃ߫��˘ā�T�?0K��$�������ˊWeL!�@b�u����T|���хI����1��ar탯{J�B��+����H����Y͙t���h�U	�oŨV�*�0��YM
����S˥Bw`��~�-4PUq]z�@)�7s�S`�p!�,c�Ѩ�c=�+�y��P��Wa���i�@lxj>��)ej�}x�7hQ�lNP��qQ��R��y�%�Tp��Nvs�m���bV@�i�<U�L�][O�'J�RM�����),��5ǅA9��*���ٚ�>U^5�����O�I,�5A�����1�#F�����n���:�@�t�tIfF����31;�9�0M�_�:,Z��v�n��_ �wHXn��	Y�%�0e4�-gݖ��4�A�ᾆ�ؤ�M�9��dr�w�����}��-򺹽�s���{`���V�7ּ:�l~J%:�C�4��bkdf���ݜ.���s�u6LH
��`���[�J�/�<J��Q�ĝt���ts�{��t'$�tF�ӛ'/ɢ�v����~")�:���� ��j�)@YʵoC-������~]硍�!���~k�	-��\��yBi�� �i��N�k�d�@�d�����Zݑ�0�4�Hb�zOt�͕GY(c�e�SML�I����K[���{m|�ۀ(n+F�`�Ԅ��H=�*���b��3�
ܧ{����֧WA���e.�I�ra��p_��i�s=���"Ƙ��&�N���`� ��.���n\��ӹp�kQ���e3R��~�8�df���mo�Yi��YC���垐#e,/o~s`�� ��+f]������	�h�?����!��\S�����<�y�^�=�n�ӑUo4k��D�)���S܎�Ro��oH/�7��~�������[��W��u`�R��~f���k40�ţ&���I��j/���ANB�٘��R�e�~	m5��^���:���r��0xx�^�-DS��	�ۥ�%i]�y����9������Gz|��RX�&������i'Q�׾�Y]g�V9�H\�6ZB:�^���֛J������t��ц3��ym��/���,0���fG�����J[�j�����1��Fg�l�=���)U-dQ3�A� ^K�#�� =�mU4_Q���Q*Q}o�kc�,Q,���R�}y&T���|�Y��G?)�n�j���%c�mW�}�����Y�?�'����L前Oe�G�"6�a����H{|���^]z�I���XK�v��9�f�t�Y�o ]��_D��������\����9�F�U0!�`2���V��_�������.3��Ҡ��C���G�^����ځ������F��+)��Y�<0 �,�5�W#x�з1
R�i3��/��W-N@NB���(m"ngH��rn5����tτN�.vƶ����s^0�7�W�d�Z���x��I�[�@�"�1�qm#�d-b�az~��=I&$6����1�{�'�s�dx|����T7|!~���T���{��}�dK�J���c�� q"������cd�[�!]57jt蓠�n(X]�ˉ��ل��t�������U$7YH����*(~(�Y�,���a�8�>��މB\X|�:F���K��zbQ���_s%5� �ԁ�|�2��Z�#e�O�j�D3�9'�j�[�|`�Vy�]����ϔ_��5�"�IVob��`'��&b�|�eE�^Ԯ�瘝D㼄n�s�/|L������z������� ��a��
�4KIa��3�0��q���9���m�:�6��~��K	}��ʒ���{#X	+;��R�@h�ϓɂ�{���o��2˗s<��t��_023��O�৞�9���(�ҜSP	 �G)Vq��	HE�ޔ �����{��6�Y������{�d��y��g�缌�򯙭 ��5K.�#L�.
Wd��D��XZçf�]���̕��Bpy]%�YQ�"Kg��b.���L�u�nΎ-]!SU](��!5�i�\��+�/��Z��FN�ʌ�`��n©�|�3'V@��y��m�G����밆螀�f�����Ƣ��5 %K����)U`ԋ��2QԢ��PTk��Fa-����f�I�=���#P5�O�"�ܘ�?��Z��j����Dtn�d�!gv�$����� �F�AC���.-��6o- sM�*���\ݚ�X�l�c�����)+�f�F���)b"����>�e����K���v��H"`kC�����57~���&�r�B�Y-H��0�Oί��l(º�?:I�$��V�[D�iL��]�zK_��m~`�T9�%VW�/|�XNx0,%�Jb����^��Wd	ء��f��m;����?�"��|ZU��R���'����\>bk�uQ ���)+R�"�:��]���?�@���.
�]�L�$�X���[/�����FK'�pn�����I4\�N�k��9W.��K����`�j�2N�̩��-�Rւl����N�I-为�ǁ����̸����V� L�ꀔJ^t58�D,;�9HY}b�R��9�=[c������N�so�ZC�&��-@w��,QC$f4a�;��&A�m%!��nW�L�m�Y��~�<3}`k$����L��S�}��|gS6�����K�R@Z�D]<<�\H�y׮]v0_�m�U�P� `R�BƄQ���?��'1jm���#2n�@����@�_��<�=����!�����"�/�u�$&x����SV�,J�=��
*j�;mF����BL$«�;�J"v�n���S�����1�h�1��r{��0��AII��-�,���Yz=/��W�-�,��;,�f�*�Ԧp����[�c\��Ȝ ٩b�T"� N��8��p����!�s���~iC"����f���&%��m����R�O�_�5~��_,%o~3��Et��6s&�mY
�L�#bn��ρ�O+]��Z�8�)���};��6���f�)��H���/x#��;9:8Ǟ2���E�I�����ր��?��%�E�?�[��>P{��/��W�R��,��'�F���zg�����5��~��$E�#;��9��΋��Mw@x'v�������ѳ�u�R�~s훫hG��U�ag7�x�c	�:b�]�i�_��}'2�\���P�`��O������.]E�XW��wߡ����HE`�!�ѱXvw{��~���k��w@
�,U� ����_��$f�ӆ_&&���ݠ�A/���M�����"�rY���[�R�	�6z0�{b��,��"I�Q�"�7�ՈҘ�_	Ŧ�/E@����O��5 '�����U
��c��k�Șk�����$��W@H�m!��qN8��ߐ�km_N�r�(� ���5�C4|ڔT9X�h�5o��{�C����ah�p�F�F�L�?w�����	����ŵ�C��d:��	,܆��+_�nm��깱EsWen�a#2{�o�.#sb��%V;Y��B�:?)p���{݆?T�/~�:ǋ9��;^3q߶2j�ۤ��G��XA=��y2�p�E$3���ύk��|W?�����gYP��;� �%P���G힢�6�_���+�&K�%�����5l�Q����{�E+/���9l���.�\��̂a��1<�6;פ������PN���+'�YPW�Ɵ��Qd]�=��W�A��^K���"2`uI �J�A>�p�JW�%����c��̍�W�#�nJ:ǶY@�l���>���*Zl���� k�w��2�n�/p^�x�Ri{�5}��0xx�F�`�N�
��c�����5"�F�ɐ���P��^�>�-����Iλ
H=Ǌ�7D�� n��:��ZlP3I:18���m�V�ѱ�X�I�o��W�	{�1x��nO�4ex�_�Z�����2D�@� /��h�2er~�@[ 2���e�J&���B tc��	+���uz�P�-]6��;tx�ى�SGP���k��Wt�sｺ��>�ނ�g�{8Pk��+5�y�jS�̋e�v�tb@�W<��Nh�<4]�L��
7H�+Y�AN ��,�i��+�t�4�1�Uv(���u��Oy��{��LXk�4L����d�>�%��*��P�z�b`��1_������u�_�y��������K$�����n��A%��<��r��tJ��L}�OH	�~1>`�>�	�+2Y�131zs�\bzN@��cL?�a�b������3�*WU7�8�*�o's�A5V3�>�s���q��?����M'�V���a�|m�gP4��K�~h�a2���>`?^@��
�B��tG��?�"�d�v�_l�;9�MO���N�ى�)������Ȱ9 {x������,zk|(��u�b��/�7��4d6�aܻZ(����<~lML8'!�C��y���nY��$�B�Ha�V�����^j��`n��&�3�s�}ß<��g��<��ˈ�	j�X�*}�"�
��@"��a��f���Q�/-�uqX���z��D`����kxACI,�����F8q(z̝x,�2(T$J�i=h6
ڜ�kuZ�ֆ)�85_7닢�֨����94��L4���
kQ��
����(Ӳ'/;ޛR6����E ��	S�:���;U��uA6^{$qn3Lt�� G��8���g��+�k+����W�w������܃�� �Y�IHQ/7�G�7�؏8�	YU�@�ߕ؋d9�g}�5�:3*ք;R[�D�u���꿜."]�����KA'����ϨX���ª52���%��Y3����4h<B�' hڸ'�3-]&�lA�u��X����z��<���%�TU�W��:n:�H����ǔ׬υ.*����'}��9H=��#�qĘ�#233�y��[���������o���5�x���
�nBc�n3��I�����׊�h���hS�c�W��-�a ����'W~ͦ1n8�%3}��S
�G�t�K}%>�^`3�B����&-��X�%� |���c�G,G���h�~�<R�Q��M�\Q��K^?o�K~*���N�Y�Փ�����2�9�?�3`��c�iG��_|q���e�A7�7����5��t������k�>߿�}+���G�=cd�qf�ɕ�~~�r0���b�	������t��#OZ��X8��{۵;{�sZ����yET\t~����*�ZX=.�~B�KiW��Dg\��/�� *$���I�1�aT�(�Eo��G�3�X���F��ײEU�3�o�um�o���X1Z�~}<x�F����7��c�5З;L��^���0گ��E�~����C�z�E�{*����[K5�uE	
�co88��'�p�rq��KF+SY����?I��w�~1�V 8�v	���åaF�E�7Kf���]���{(ģx�ڎ�����x&пbG����XY뢢J�S�4i���ג�tǱT�Vj�h�^��BU��L�~@�Z�or|�y��@�z IAܒ�x���>��y!K��1�clF��am$O�ۮ�u�.Q!�U�l���F��R��kh��� !�t���r!���4�
���^$P�ds��P�u;�9��_�pA��>)���~b_��C�@o�O��P�[�Eo�VhK���<�5������_��G���nɤ��{��̡Rz�u��f0�8�RD�S 5{�:53{&���m�2�F�{���,��i��-t*v.ǯ�
E�Tu�Uk��(�4��a�I�R���~�P��|��=z��_��FV�5P`$��+4~���1��k/���u(�@�Ϊ�Hv����Q��Vl�A�l�}��K� ����@��|�y��]\Ƒ����B2��+M0!H%��+��\����\��tX�K�t������?5BVyX�f|��$��(s�2e���o�����C8E����ⷌ�L}`'1g ����ԁ�Y-��i���BK�r0�;FX]���_�Z"�ɗ��X�Uc�)7-`�K�����ֳ�߲7����q�P9�N�4�b�2�k���ױ��������Q�y���A�����Ѹ���Xjd@�R�C�q��jݢ`T$��fe�s�G��4u�o��(����´<��aW+��"@�p�`)����f�	c d5�r]Έ���o�:�R�`�x�U_:擾t�?�RG���%h7X�E�Y���<A��V�;Y��KVZ֧x��3u�+���:�lIQ��3�|�G��
�=��&J��Ӯ-x:��^wx��݂���C�C��)��Kt5V����Ez��n�*ǯ���"��M�M�W���<be����-�i���qK�V��y�2O«���u���6�r*��Ҽ�\����ڱ+�nG�c���.9O�B���y��!�Н��k��q|�
�`�:�	uW�2����6Vt+��~f���p]0Z�%�M�ۑ{.ʌb�%�?֧��
2{�,�+ �~7��Vl_$v�֘;���ҙm-��7�ƈя|�K�}!�^˫�B��@׆0�b[x��t�[`��4FOx��/� �}��=�B�5C,o1�{�rӵ�3#~#�1�?���Q7��AĮ�X$�T�m��Z�`"A����e�S�f����2H�L�ÝS��H��G�N��	�c�e[���Zs����O)�L����#CW��[�v���b�T[u@����, @����RŘs4�/������Z�z�	Z�d�yk_?-l���z��&�o��U��f��Y��	̡��T�*/��G�f���+�0�/3�y���:����AxX�?U�X�9�N�	$�֤��h \�2U�Z�I�eA��+B�TG[�"i�* I�����H���.j�Q��H���]\Jz01����}���N$&����z�]4j����w�W?�! ���W�+��N�,����\������RD�&])��/D�F�����j�a�ZO���枈2�E�asMt+?� k���ji����T�x8��@kK��S�?G�a8��7c��Lc�����\��Ȕ�
,h��@uF9�e+�+'�d舖�u����V��nS�D��[t[�5MIԭ�z��Y@WZ�$a���I�0��:���{n7�,��5* y:�"]����8�oRPpw���`w*{๡���e:Ѥ=��������Qy�&f	��Z1�E�H��?]BS�:2�� �"��t�+M���0^���p̥�Ųb&���0�M��'��܃̅V�Tt6��0B_��ΐ᳉J�����T�Q�b�
Ѿ?��6M!0���2��tb��(�nE�c?�m����֔D`�[��^�l�z���攴d�0�c��!jf���ǽ�32�WKO؁�@C�2pڬ6�BX�и�7?7���N]-J�\�řg.��E��^}T0�@3=�B���s��kV�gXf�W�N��O����n���p��WTI&;2���ޜ�I;:�;����UnD�C;K�p�f�Vzm�r��K�ӟ��}c��O��*��dJ����)lLj��c�b��k��㮂Y�R-۱&V�ݑ�bR�'����$0������7+�1��`����bǀ�4E���v����G|�P�ܯ�9M��)�c�Ą����Abx�=�fD�7� ���gƂ�xz�J�݉��r�*�:;;��=�ǱWa9�@`�W�='�=f4d>�\{�\����1��(�:먪�ƍ+u	tD��tg��"#�B�w3*fB`D���-��O+���=��7���~���v�77f[�u |�/�%~؇�w���y�X$1��g�#�"�
��G�&���S���O� �hڊ((Q���T&!+��Й]�Z�ڙcDf ��8�hJ���ݛb5zh�hmZ��[�[g�߸�E���P��!Q]1�5�V�~���*��ۺ`��P��u�*[�+
����;i�6�sЀ��#4.�AB�+�l��Y�z��}��,`�~�I
J2�W�|�)�>5W7гsaʖh}h�%m��%tư�/½���01ȁ`~g�(岦y��������0ϱ�8��ZO�7b�G�L C>���3��N ��6��"������>B�@;x�=p���ş�tb�ɪ�yye�����*ȧ���\�35��?2ުfW�D��4�CFz��vt���^�����2��"T�5��
˂�8�"�j`s��v��7L5)��5�<�e���r5�k��������r�1+g��_���5�V��+�"��ӆ&�t���uK��Q�>
��y�������9���I��D�*@ǅ�0�=��*(�U(�{�F(ݵ��ˌH�=����hgqN���(s==���������4��\XZ���;)��|^z�5��ۗ�`/�K/��E���*ZW'�C\Dw�h@{`�es���A�/��3�y �Ź2�t��[���5>\�"�q����ٹ(��G�CY�A�4X�@�
���7�H�&���E�H~$��B�̵U�k>)�oO݅�����:�7��o�Ű�����}��ol}��ZJ���V��b�J�G�p.��F�Ӝ4�3�C���gy�
����!l�KQ6�-#7 �,W=�����A���췸�0��Y ��
K��F,���՟�������:Y�ΊUeja������=��Z��k��� �9�2x3��Y��j���2�&�xj�����W09�L�M'�r�jpC�����I`j�X(bN8��v�R��5�л����ҿ����w���JA����1�x���(H/RҞ���Ex1��7�G �*�Ot,��H���Y\�Ӊ!0�e��{���ļ����O�2s�d�%^ΪcD5��{��&�xu�E���k���lJV������}�"�
����E�#
͠�z<u �ʯ���Ѧ�����<+��!�X+���B��Y�
۔���	�Ko��(Q7x;,2��T0��c��/\���A�2�)�,��X0�A���/  S�f�*�������M]�������u�.��.Q����]��q��1��:�T��dʆ̀� �@�!a�ہP���w��Y�ۻ�g|�U vI<�W�lV�s��׀3�p�b�\IMך؟k7�>��f�B�T�'���j�7L�<ˠm@$�h�������c�#�g��m�Z��N�o��}�%���y���xa8���r��]m�.��M$ˈ��/�`�(���	�eKש�ϕ4@��\���8��F��:��"���u�����F��%�ei��ޗ��sR����a.��s��a]U��+.P@X���&���!�C��jB^`����I�d-�P
��O#V��,�t��w|�Q>�=.]�S�ص��%��Ӭ��v�q�������`r�M��)���<.�hlN/�#{`�JG-�A)9Ī1%��]��І(	:I�˰�Bvd�0�0��;�κN	��0-�M��3O�����@�����$��:����-�� P����P��K��h���^K:�A
�C�@1:�R*�fR?��v=�z�:���6�q9�_��͵Ⱦ��(�^��.U�d���� �im�!&�ĭG���\��OXA��S����9�o��a{|�j�g-�ݴ�Į	���Wg�#����e�w��vG끅�1_���j�X��V}�R�^|"Ѕ�����F��Kc��˗C}�0����G����ʌ�b�U�0>�j�\���NO�˜���c6-�:�6#�)��I��xr/S�n�|��V�=�o�����?��|=R1ٙ���n�U8���%T�eK�ʆ�;�~s�~��Ɯ�U������Q�JF��⩣��W)_1=�j'4�
\�����@#efgU�@��b�5b 	�+']?��~,�i���X >:�k�ʫφ)K�43�؝kg1�R��&�������<�SW�;�@,s�	ۭ�]�ELW��]|�ؗֈ�������O�TL(ሻn+�"����v�~z?��̛=	rF�R��K8pC��G�N�aQ��Q�d:���H4��SK��ۧ��g���F���	���0�������.�[TW�ɻ��ɷ}ձJ��Ho142�4��ѻI ��W��->��Q~��J2�F�Kx�Y�ƚ�R9S27��}��v��L/]�࢞K?y�rB܉���Q�3��p:{��% /��fϤs��W�>|Iޒ��.���Xu��~�DfK$ 0���X�c��qP5�[��ދc`N�p��bB�C���*fּa����dw�)L_��&�m|q!�}�¤T��\A���Nf���dr�;e�d��7�4MT.��Yl��]�^0W)aW���;�=w�Z����()�XJ׍����+~u��N
�9�MkaǹM�Ǿ������ڞy{b{b�r�&l��|���h@ޗ���������0����
�O|���XR��؊Џ��������,6��ƾ4J|�ޑM1�fU�ǚ��b�FYۧp��_�&��ˬE!�B��/������mǩ��u  ��غ��|�T��q)s�z7��\i^'��U_C�ٔ��7m���I}�=��a1VB�1��j_p]܀Q���{��$�/DF�G�l�k�.��Ȗʦ�t��R��\\59�/3���'����R�b��}kDrC(�b�H�i���U/+��Q�:,$��+��?��m�(�of�����_،޷�~C[��^��ֽ�m�Ro0I���G�L���Ru�����G�ؙ��tg	��&��,��%�z�;�.��tE9�	}(����t��P��� G}jjY�(�'��n��V|7�bۃ�|%��O�`��޾�-*�=Z�=2�ݠO��������������j�@'x�4����A�%�	�b�2���G������w_Y���Mw1���ݷ$)�@��  ��ЏM�76����K�\q1p���Ll<b���Te��R |sp�_'�=pg��9����`�,������~���� �)�'a��>�bC�!f�A��܊a]�8�=�7 �z/��L��A�B=b?��琱�'�
"��G�!~��)�j��)k�}���y3Ԫ�0�%�ǞS!��wX[8�a\G֋ǀA|A�*r�����}F+m�Е�Gr{r�
S�MV|��G"`%�J-)fo�bu�����][f�8>�_DG$ �r�3eZ���2l��G��aD*�f�Y��Y�"&���eH�?7�ss��h��J��v5�b�Z�O�F�:Z:o\�8p�ފ�����Ksĕw|�,����"�&� W�vo����)�)#��Q
����ш����sXU�ʖM IQ!¯R�Z7t��������Q!��P2Z��~���]=��ÀY��{�`��b��K[��R<���I����&MQ^_��j���0��kQ�RK�1>���
S�~*�� �[���0�=
ZƼLR����9*PY;�~����E`���<�����qV؃Y�~�_ n��z�>P�5
���Kѥ`1��-̸���|��
���#��OU$D7�L�+�d��9��N�^�B���d�i)l�d��p�����O���]���3�t��ġ���(io�N�E�#2R
�)uD[b�I�m'0	��]O1��u����~S}1>;���wR%X�`�C1�A�Z�\���vHFD���?y�)�J�!dkt�5nt󭋨�����w����0U���LqZ����df7Mw�?Ǖ�����^��ӫ0�Ӝ�����W$.G�v�4Z���A%y_�_��;h�.G��c�M�/����hJN�4�p����)��;{ h�s�@��K�����h��A=�J�|#?zib�رl��.�������~��6oƮ��r��ߣ�OD�0+fg����K`s���L1X���<Ĵlk�N��z�)ۢ�:8J��}��K�v +�;JXh&)3=��4�̂D�C�*�ЬCpgaK(�U()lW�X��hq�+:AN`-�]v����Ǯ�Iht�Q!��:ox5�/���,��ϴ�X�Z��Y� �_x�e�%w��O����oa�I+�e���G{�̶�:� #sR�>o��N���/����߹��F`4	ˉ�y���k���}��M��ypX�[<t�B�^�����0�!���p�B�ۤϋ8���ߍ���8q$J�3��DU��5��A��=u��ya;Һ�>�<�xإ���~v���ۖ<ԉN��6�ҏ�.F#
@]�d.�PB����p@uh��<���܏`k�2���SvV�� ��2�����&I	�=ϴ��t9Fݮj}K��D�|u$a�m����$λ�K�"�A����10���5���W��;{Q�LΒw6�Ѝ�h��u�Tc6���$�0�$�K8N�2��}�d�}��w�i�'S�^❩I�Ym���0d�)��Y�E y0�<ZjY��{;���$M��xX���{nU���<��@��4B�i�{��ߤVX�7]�4�_�:P����Ki��B�k���an�=�������8�K��\�1Pt��Ž��T��9��#��I�����K\�k��ʩfq��Q�K%��vv��q/���� � �@��v��t��ZE��d,@�0wZ�����<ge7��+\�F7|�E�3}y�����T�,���jn��٣�0���z�ɪ�~��dyW�k���m���(>�R:y��&8m�,Fq�&���_��@���U1��J�_�?�����	�9E�Ϯ����)��׳��`'�i/E�@n#�47s�Y;��.���R*�f��CXs���f$瓷 c�@M��YbS����7;�:���K`!a		J�ak��$T�u�>�ĉ0�d�޷r�����K��=��.���oL�>��@�������AU�	p�T��;��I,����G���x�.���%;1�5S�� -$:H�?�s'V������&&f�=k�$
��ֻL�4�:���*ҡ�F ��<���lS�sM���1���3Ӗ�l�����S';�_>������J���_(]�:ꜧ@W� 31c�q��v�M�Rn�]�ƚd��d<p|���SB�X�sL�<>la��-�p�;�b�� I��g9L�~��Ί%׹-��@�N�h�M�l��Q\g{�H�ߞgJ��5ƞ�1\��Ii�T;@�⌸���A��-e�Q�����_�&�Y%�N�˿^�,��?/>26�=w\�����1T��O��JV�����1��,���)��:T�����O	���</�l3��+���a`��`f�no<f� �	[`)P�n�iȻ�0��4K}��� �l���������0�n�m*$\����SJ��o�o	7-��\�J�.�+�6� G�-_h��Y9^��5G�Si��O$�*���u33�?X�@̧J,+~�{>P%J*l��H��K��(Nw���8��An~�y�|ՠ�dIr�XȦ�1�������4�~{V�~�QɕN�.ě��2��b�����l�.;��(�P6��%l��� t��Ϻ�jr#��wͧp@�� ��jDf�����t=�ٜ,�m��u�L��o�C�6�u�)�C"N�d\�i������JV�F:< DF��DZM6�^�9��}���Xb�m�ֽ*#��3t�a��������>:z�}�� -v,�x1��!8��3_��cǯ��.e��W�#�J�n�DxC�+��Jʍ��,����i��$eYU<u"^��ɳ�X�Ǒ��؏�r"/���D	
�vԈ�X7�Y.H4k�r���(`V��
�ʐԴ�	R��WSv-�S��{�z��/!��۫[�[2�e����X۶�/���(�Z\�z�繠h ��L��4��6N�-��D��J����;C���hټ�_�Y��|;\��
�������0ٲ�=���� �D�8��X��8C���8���7M�@�y�6Vb����4�Y���߈,WO.�'Ӫ_�eUb{3����[:�ҕ�y��.��oL[Þ�P�q�f�oݽZu���r#���ɞ�9)�!�v/D-�	�������yD tpf=�^����t��xC)�dO�Β�x�f㱆��v�e��e���	�~
���A��#/-�SB�Ɍ�^�x�{	�C$Gg"�_�t qR�O5����Q�)�Ug8��=<I��b|6h���b�Ԩ����	������'�n�r�ݶX���r�ۅ�%'�w�J
��9�H���1*2�/��''��ktDy�Z�~7��86��d/�^�!�P���Sǰ39v���s�H�	�� $�������C*����}G;���Zu��=��S��4�U?�̤����$vce�5�ȒG���L�����<�5?3t��A����TR<�숌T�g(�?�����;z�5���7�� &���a�-؆�pz�q=F�� o�=��s��aA�o
;��f#"��0�qd,+��Kw�5���G�1T���1$�~E�B̭�6M�
k�|������-�Q�E7)V���}���T�����Tٱ��&d���
S�V���G��U��
-�{�gz[%�&��)K�su�O�j>���<����	���$������$�����Vz ��<��Ǌ��>��}��쑅*։Jv�bc�~�4���^����g�2-ea�*�vzu�M��% �>\��V���
�Q��܇P:�lh^�=���_��*0�h�*�[�c�|�E0�#0}u��D_Q���Ye�"4���@��{�L@4d���*Aa�q�3>&��>άI�����2qr��=9�!�����g��������W`z���n��W���ܳ�T����PWfEtAP�2��y�ͺ`��F&�T-�*�?���������{iN*�w��⊲tÐ:���/�cNe��EB��N�,��K��8�cg�/U�ϣ��uk�4��%`e7|"ޭ��}����u5:��w/�>=�.P:WLN�N��`�>sJ�dD�Vi=XDvS(�Z]��|'9��\�,P�� ����Q&�л�(�5,������"tM��� ��Q�y�/v4��sy��lF��O��Ud �د峀5��@J��ڥ���8es@=_��ؘ	A@	���9�-!�U�U��DA1�o6S-?�h�M0(��n�-1��j3t�ތ�\���V������Ɔ������3��u\`	��#�������E����foI	,���M�/�m̟�#M0�%o�<�l}z*nR�њ2�\z�3m�ue�dX��6�K�E����| SaI���]F���3�Я N'y����9�
����Ǿ�p~�R�;��>953�;�I���dE�x_�P� �]N�T�������ʂ�M�X_�k�}���C����_�{0�h{6�R�%������4�(ᕜ��{�� ���}��%bh�$���ұg�_d����Gz}�xo�sq����(�{��f
�^�Ζm4(�I����������A�QI_}>�"��E�s�Y-�ǠI@6�[kwʻfaJ6����=�X%20!u�e�� ߑL��3I��5�D�-�X~:�n����Z*VT����j�@/�{0
Q ��3M�m~X�3�z��͍�E�_�� I6|������)�n��Č-B(��4����]���b��?��_����I����J�2쟲��}2n�A�>51&-��CP��p�����a`�K ��� n��"��?�`W�������x��_�G7e�	����<���x��n��)�OZ�ᶔ:��/1C���Z����*�k���/؈�d޺��R���X�[ʺ�Mh���%Α3�e*+Ǉ�<I>�0nz���:��[�0#I�[��?��7W��Z��(�w��P���b�tب���&���s*Dx0{�n|@�[U�V�Z�R���gvN�$%� ҙ�1$M��8���2]y셏K.qp8Z]�gMpPݵ^���89E�K�ZQ�h0�_)�:uJi�|�s�*ƈTc^��"�,}(K�^h#���ޭ�p+3my�I
��}�ZG�S���9?�Cx_��xE?��(y%�EoHe�R�P�BKA�o�yοO$�}�͝Buc8JK ���!ľ.Ҕ��֖	Ep߾r�%����[U�;A�yH�Z�{7�_󋾾��+��=��^���.^{1����b��{����R��tcH*��R�/Ѵ�'���|���opJ����3Gp�r�+�E&������� ���/�j`T�9��C�26<��Y=-gL�i����!�b�����C��DTɧ�`�8WW!%�P������,�/�X����$��%*c�m��W ����>=��1J��ij��y݌O��%���bTϚO�ô������Zأ����it���tq�������i�GhK�TU<sa�`~,�}��8����m�o���ā����\-��L�6$=W����)�0��V`��&��8��&�(�	�Ɲ+�����"���)��B�ϡ� �4�{�A�',u֔�qc�@զ@��:3��5�k�f�,��1�L_�5�DQ�ᪧ�f96� �w����uΈ�u\�'��ߴ�<�Q]܇ZX!ʤv~����Q����A^�aa�U;�MH=`��0ӻ�m�AI�&��T�AZͅЛZ6<s.U���=�1L�aaVZ����Lz�����9�B��H� mN�rnά�F.�sI��<E�� �Z����5��gR�oL������#B/⶯GT7b,l$c\?j����N3ov�y<���K�۱�ۛ��TX������n�:���ר"9)���t7�o��=�u��z��}4�_P{j�N,W�Sg�LL?!�C:� � IW�v�o��t��e^L���a��e���C����hp��SN%��PP��u͓�죄T�%�䯐~���p�`V�G�CJ������=ς�@�j�	����M9?~_�#k�G�>���H�w -H�G?O�[����?%�Y�笣��?k�5�~�d��]F�Т/ӽU/+������jk^�n	H[@ߛ��7����@ro�9S5ecJR �[�Vx��j����e���\�2��lTA��ߑ��S���p���>��cU��kw����P����eXf��6{	G�/Wd�SF���|�%�;'C��S�R�f6����x��,JA�~*^4�EVr�v�h�����������Q)�RjM5'���\�U�z�� ��$��iq`
f3w׈�m�n�]W`��,��.���~�(�?0�b�ы��Ø�l�
z,Sht.{�$�����f�	���|9��.5���F�ҖL�p«S-�����q���w|S齎���w�exL��J�Q`�� �[��l1@�pTr�"Z)�'{��_�X9��o���B>�q1At�?�,EݧF�%f�K{x����o�M�G��ӎDK���a<N�y�;����1<�^�3U���.�%9��=h��Ӥ�Z�]֩���R|�Y]������I!�`���"�E�-��Uw�=�5��F�	G,WD'[R�,A���|�ފd�f6][�^q������'����Y)-��ڂO�}�6���0����lG��n�b����6q+����*:j��+�CT�A�K�&G�hJn\�|k�%O��`k&��Y��]�/Sʺ2y��T/3!�L�����C�踩p@ν���J%���bpQ0�'W���[��,��A�H`�>c����p�9r(��{lM���"K-�6��+E�̙ݠ'q�R�ހ��wӲxV�0�&V�a�YŨzw5�g�8m~���On\����!bW+�:}q��]��흓Þ���?lI�l�|�PuG{�����h��7�,2���]dȾˍ�@�L��o�M��[�o�R�;���:�J�����}�2���3�Ȃ��]�v-�_��Hx�I?�ᾊ���Td[_�l7���H�1��d�nO�Px�j�ףqZ�����t�e����($"��-�>������Oqf,쿓�Ŀ����jَ�[�֬�͏	�Q��v]�⎼ne���M���M;�RQv$R�e�Ä�����Լ�2#�,�����M�cߵK�0���ͣ(���N�d�8%�Ԍ����.�$~M�Up��SHz��`7f��G�����9>��������f��-Ew^���ĉ7����.TT�_�Ҍa?�!ә�a"���9уs�G�m���yé�e�ձb��r/H���+��W��I'6$�0��i�_�9I�n'~�z�;}�է����~��^˻v������e�iN����c�����Bd*�T?���OA��aɡ�_�T&�ML��婸G���sv����r���̶��E��QD�Q�t��d��Z�z�^!,�1���e9Ξ��֯6ܧ ��~=@��Ph�#��3Q��F��N]�?i�<J��c;��ߩJ�@D4k=
`�|���F�(���|}��޼�^��<�m?���Q{����H�{Xx���I�	k��װ[W?�NUx�f�ȹ�g�ȃ��|t��|�yA�G����;���.�����L]g@SK�zp�WT�#]����H�%@�*R�HU��T��� ���*]BQB�Є�B�s�����_����g�yf��l�5�ʟU�����&IN�Ck�����~r�}EkĎ?/n�SU�����荗����X��7���[w"p���JzL;�^�"���ފ�j��`I�;��z���R����(S[Hș�Wӱv�xq��*K:k���#�1/ialU?���3����	���C\�d�򡶹>��\I5Ë:��Zx�bП�x-�#C�τE��:�E;A��A��!*��Rj��2��H%��/���,���%M�f&�:g?�,�B�F�CD�1Ĳ��oNm���h=Gm��f�Xv���S�0�Deݭ��P5��.�ZC���0�5���ӟW�pդ��E`���\�`�+����[�_L�/W��s4�u�p%�tj���ꃡ��<�aL�L�8m�����������<���Ǔ��,�¡չ=К>�(շ$�����F'�<CG����`ӛ��_�����|��%���ak0�X&6|�a��ҀxQc�𔲋�/d\�j�S�K#)h%�le��[-8��s;�^`%���9D���w�hzuJvP��UX���vJ���{j����w�{��?���,���w?�ΆPY���w�[ pgW/�F�à�&|��c�h��{�J�*N2q�JR}p��OwkON�S�����|%�c�_9�5�ܘ��-�㿙7q�H�L�G:���'U1i�C�x<�Y�����i��n���w� ��V�z�Q0j�����9�����C���Y�z"4D1Kv�x�8�b:�;Ow"o=�ey�ѬL����2���������v�,��q5W0G"��,�c�,H~���Y�=c��^������Z��Y�ŽmG�[�IX*�y+����N�k�2E�2C	R���b�������"BjI��+P��O��v�d��F[�����/�Q�N6�BO(���p�j�q����TNI�De{|��]�q�	����_dw��/����[��m����d.������d���W�G��
�� Ȼ�k��/��Rv��~�����p�1����PA��'O�Y���`�Ef��ӧ��^��3�^����ͲK�oM�@5��im%4�C��٫0��T?W!()	j,iF`:�dW��aQ/���k�S���R�����S�/�:Q��z�~��_ӘO��hN�B����w�臒/�3(��%�]���}������l�;S����6�#��OR�2���)Kfd$�[����Ǝ�M8��)Rᡄ?�*[L�$'�tL�-��d���$�oX  =��w��7���Y���jK��qP{�s��h�R�ehȍ�w�q 	ժ1ۅ���rL�.o:�դ)[*�P��QO%�`��O��HH �F�ͤe5�Q�p/���b3	���EHL�#n�{.��FD�do۹?�j�����<$2�CO���kE*�~�����Y��Crá���/M�k�gቢ��/:ܥ��82�I=q�ܨ�#���my��Q�~S�\2(��`:��p� �wH����UR��j�nOB�CO5��[K�\5}��6^�ýt��Gv2U�=��rM��mԺ��K��ˎ�rF_|��Jz��bה�,ڹI��ڷEY8s��˗]̤w>�b�@��r�H/j�iLY������&�r������l�ܝH1n�R�~;
״���KL�Qo]e�[TVx���Z�3�l�V�����2U�
��g����I���:�w�4ńN���;*��.1�>4��{�LLf�잦|��7�|8ו�*��X�qys����F<�n��@A�M�0g����p���j��c��֛�N��}�'
y!r��ñ�x�4a�RH���5�<���kQ�i��]a;�ұ�ר�zxv���G��\���0�J5�!��Gn1\[�{Wlne� �ֈ63力������:�j�A��,��nZ4��:B��!��~�s��E6��~���k9���q���)�uAuQ�Bߴ�w��s�}�'�'���1S\�����t�s×r���IGs�!?�o��n_Mk��l$<�YX#q��F,��V'�gT�O'3������홚S'��u�:�o[xڂ�֪�nb��+$3������G/��y_3�|a�[TS��^͕l�<m ګ�Ng݅�-��b��ܧ�aGX+B|�``��dm4��^p�.b�o��B��S5��B=��C�4�J~�_ۚ�",���th����]�$�v��c���n�P8d��?7���`��r	�R[�;E*f�M�F�R���e�M�����K�\j����/�����9 ��)h���r��T�����.$�4�nLn��¹�����*1��?����s��e��{eQ��S��l�����|����,!�:�{�~o!�J�e�Ulg�FV�>Io��0�W3��9Xp���ҽ�m����(�^&E]��-�*�{���4��nǔJ1S���
6����8΃�߇B|B��T~�@_D�a%o�������exa�����.D|�(�r��Q	�~���~�z��0������@�?T̀�t��i�.��x�2,)����q�6�~V��:�g�S�+�J`U����������B��I��Q�;/�wj	����*� ��̝�.�f�c���'����졧����K=��/���'~�͝:ع�͌������Oy��8�����H�!)|�{�uS���$�t;-�:����.�X?�=�,^Xmdˏ"�=���y���j<G���A0�<��d8����������#��MUbp� �irgP�Wv&���_�Ty{����Ub�a Csc�
�mK�F�"������lV�(���X?���f�e�j]#�c�}a�k`3� S��%��T{7��z{������j;)��&�[u@�ؘA���܏ˑu5R���<-}� l߻��(^�tW6�&,�*����{��R�ù��g�����&�k�Hy%y@v9S׹�+�X��]!�rݗ"�Dn�ٔ,尞��.�T�v�j���9f� R-{�폿F����"���h�rs��5��{�$��6{��🙏�<>z���i���&7g������z���$�2z�V�a\�i�_"����^�D��!�=p$#Ƽ#�Y�5�;�ʥu�DR���3��\y�Nuk"��J���ߔ�b]��	������� U�:�ͺ� �OR�FKLב�2�{(S��)���,�6��4�Epq2Q�����ґM��&yl]� �9�F�a�ȥ���8�d����>�:���=�9�5��R�nkF&�i竷?b(�4n�IM����FU&��'��Jz��E�{ y�6���7�L~��[d�0'��tXVb`���(���Q8/�����K�Y���b��6J��6a�C�в.aN0l(����0��F$%��)w��4A�C!"
��g�ٱQ]�j��O:ʮR��SZ���(��j��<�����M9�]m94�!rlA��U����M�YC�Ő�N�ڊR�d)�j����BOdꩄ�����y�wI�/�A?0�暆x��j)�~�F��K��r׍���w.,�P<靬��������� ���l}����#�2�u�x��;t�T�@پS�q�q����A�܁Ef��|���l�׀Ph.��h�\��F�g�۫.�r&a������-r�\X����t�0M�iD�v�@�*�|y	��]�MO8?^�H辐�6&(.\OpM��e&���0}��L9n�F�j�����Zy��(?��!iy�g*��u��]��A�H!�{�d�};L����'��_��6�|�z�#�R#�C'�ö��F��&"�+Q�&^��@�I��1P>��N���2n`0�Nh�q�8�A[Š��9,*rf#��3,C� Ȟ]UW<~������j��hZ�����)�)Z��+ǜ�����閕�����
�J- ����m�a]&&�*)��^��g.�5�S�(�uR��y=�3����Wz��Op��LR*]
�F4X	8�᡽[�Cjʳ.#�A����Jg�f�|8���m���`$���\����Մ��/@(��髊��B{�81��,eg:ږ��^ؓk�����)>½qw_qcLy�7ִ�����*�F+�_�Nz$���%P�bܡ�mQh�{�QH1L�Kr��G.;JVPP�ӻ7�d?nw����)���G쎢��:��8q[ա��@���##t�~((5��Zb���g�=�]
���:!T.ܨf|~����["e����L3_��s�=�$=E7&��m��w������4]�wvDu�Q�Qo����(wJg�a�'MS��rW|h��?���ri>!���#���U��j�k�.���x��ZW1`�9y�x?��Iʩ����yR��g���P� 
̋��5����/ov��+X�Fp���^��؀��=�T]נ����)��T��.0
v�����L�)�Jn_S�hn:S�(}���eV7�J�F�uj��;����kzG���nρ�����g#��{�pW���������("��S�n�O��r#��0�� mM��
����<g*\2�Cʪ��t���1̸RQt|p�DT�����9�.����l���2�m�{�4"C^^uN�j��� z-�mexlnC�,Ě�mM�	�2~%t@}�#T���1ԕ�� ��2%��v�>hD{��m���9����0})*���ٸEr�ۯ�_w���lqj��L`�2�#���7�����8�Zbo��!�"�lI�Q������p9�f���z�h�:�3T:^�%i���CL���V��I�f �����
 ?�V� ���ٯ��������"j�J�j�1`�+OU]�	���&��$���o� �>�r��ӫ��:T0����{�q�[!A����P�S��B_5��	�.\.x-�,��&�cQA�۩<ˏ�D�t�����x�}�;Y,��s��,�&y�_���2��`_���������0ec@����U���)��az��ś��DG����z�@?��n�ݬ� �*1c`����|���U=]����>�z$ʏ8D�O����1�L�Y��pTh�s�؞vL�z��2���Ӳ�,8������ah��z;���������rz���e�$ߧD?�z�qAXJU2�4�xSx����ԣZ[,v_�E<���A|�T �*m:^�p��B�+<�]NԵ$�E%����1fU�1!�8ꦵ RWQF�P@���['�z�{����L\�g�Pu��r�MExkOB����aJ�xi35˒�D��&%�Q>o��]����j��r�vmI���-{�tN��_i��.p�c�*IN�(v��=�K��4���{1�� ~� ���N�MNޱ��֡��,yv�o�%�<땘eQ�n��Aj���E%���:_�t[�|l������ش&�m=KrI]"�J2���v.����/B5�>�����D:�*�ѵ����cB�3��j��
-�md���F�w��SAv/�D��y`�X�BST����H{���y���G.�:z�r�Ʒ{�[q
�g<7�N8�r��V�����?_��=	��aJϺ*C_�k�J���2�O�	������N��w ������_V�ߌ3z��#Ǥ&��T{����[;�q��do��M��nRC�@���i�U���&����>k7�\pB�>���	?r#3͇'N��!�g8�S�2�+�;�h޵�M�.�1㹕z����% F���V���F��Kn��H�<�*�����.{K/jq;Jͤ�Zp��I�`�}��3�/�veZx��g�� ��XL(��	g�P}�/�?$u�KWn�x�neMyG�6���j7<��C��i�n�:TmE�y�
�"�����Y�DR~/����	쓜�7ZN���ݪ�u�_�A�+<m#	.W�*��[U���k�/#?����|E n�������P&8}ڴ���١^�T-��_�CC�'5�(�������8r.����p���0h=���"W?��九92j�Q	�`#8��j��:&4J�^]�Lv�ڮ"�^`2�}YnKy�`����j�����,3�f{�+���\�"2n�^(��}M���΢�}�ۀ��8��p����
�Qe`5m�������M�򑬲�	�K+�����%H��q�É�����,�X�K�7�lPsç�څY�
%K���K7�����r���k�5�|���������X�>s�V��m�&2i��Y�>f���j�[M�QS�����ޠ.H�ʻ��[ėԺ�c�D�2�[��F�MI�4[��G�ؤ�
e^k���'�H�)M�1h3��YL!�J~d��#���i�hu���l��GF$��|��]U�(�4h�2��ת�:����P]cW����9��3���N�QI�G�L�dW'����˛�C#���N�\v��O\�?9���_���¸FX���Ϭ%�]��g���eO�a���	YJC�Т8ز!@�Zʟ�,�HK�	>�nJ<��$������y�W�`M�HSf<���a#���gx��P�^$�~6�-(74��FI1y3Ћ�gc9������+]�-�0W0�F$wΠJ��� ����e�N���|Q��m�]�jS��$
���C����j�2����/9�G���i�z77�J3�|I��̘��KD�����*����#��d����1�c��M�6nfk��y:|�f�慽���{G���lYa¼�9����痍��e����A�nGnj���G�\YS
����r�˸���������z�|���PY��~L�,[�u�Ӎ��z��2)4���}�c�7���"#u��4(XD����W�gs��Ն��Y�渽_���T�1�(�,�M�u��n������9 #���,�����Z�3���FB���o��IĬ8�dx��e�]�ɗ�.����Ӹqw�:�j��DͷM�gHс!^rݠj��W*���RTf�G_.k�qs�P�rØ�5���W*��,�}߷��%~ ����;��u3�9yJ~^}�ߨP����1��*�%[�6d�q�ɼ88�}���l�@,p�qP��l�;L�C�Y6���������C�{9�����oR3)���v�������l�_Բ�z�6����>�Qg��;0�6*R��P$q�CTJ(�W�iŐ�>n	�#T�O�0}3ں����0�=������5:�y@�d�&P� �ƻT��)�R5䗖�r���X������U�Z�o�p�e-��z�ㄇ��J,�����N�Z$���a>�G>��?M+_a9��Ѥ��\ڼnĂ�-	�M���Ɨ�3��8��^,������v�R��f�/�W���C�F7��}Ɨ���Mi�
)�ZZC�}��(�C��eٵ*_��~�oOIs?�Q�k:��f�!��b��^�d�Y�x�AQd�2�\�	�K�1|�,<'&�IPG��{���c9�o�Nyp���pA6��國�rp}o�ދA��ܢ�-��z�;�d�*�� 8)�Ƃ\
I��[&��ܬ:3D�E�lne�i�ť�]5�18۵��L#?��6��f��t+ �E����*���"���b����?�e�!��3��v0������0���nￛ"U��X���6���l���E�h� �b��4�c�>q�R�#ұ�g��Mr�:,9K� W�(n%,P�U�ۭkO[6C��vEwx�����K�)�k�^��:�fB�D��[$hKM��m���L�d	���\��u�gX�(�Pi!�d�������T�3BnrM��4n0�n�.w�[e��c�G�긆_�Ҿ���I|�;w3��rQwb��ln��0_��@��Y�Qu�o�x����<3�����R2�aBh��X��ݖEn2���(�epdT0��(�.:�A�˲�_�}�4-��P�	[��"�R�@Y�=?ˇ���L����d��G�tϘ��B�kD�|�J�1)�]?�k���T(1�8r���͘�[_�姧Y�J��o�w��� )ȕkn����+��)Ϳ���+DV.2Ⱥ��od����I���G�o��MQ�oˢ��8��1�JJ@���==fQ�����+�\	�x��gW$}M�V�'+n��2 ��ضi_�?�j@��1;Q�e~�,�=�vX����Dc��+�!@�W�7́����]��GG�� o*�\�E��4 ^-�p��`�j��綛���g���Ik�kqN"!y*�۫������M�hXq3�������LU/y4ÂWsbb��3���""\�jo��T����<�?03�0�|�ċ޺L�q���ejw[�bej�0�f�|���mI�$s&���l-<x��Q����Q���f��\�ࢥ��^rrm�H����n�@�٣R0���U���I�?�S`Zn\/�vhls����xteed�3S�|ߺ�ұi��@,|1'\�2h�b����!n7�������O�P�ݫ�XZ�����Ր�Q�Uh��8 �[K�����WVG��ip��Y��ay˽
R�h�oX�� �Z�f��Hi�\,9� �"�Qt��9S �"�����BYt'c�ٴL"�DR<�J=�9z��P
]�/$mT��h�����w�7|=IN;�MXk�T�)ﺆ݃�f��.����7e�V���>�Z*A�l�=;ԩ�:|�=�����J�M^d��J��Zښ̴�s:=�5��p`���Ȱ�T�3�����%�O:�ԭ�o=2�o[�p��d�x�`�)]L�<G��	(R���v���)p];��4�4j)L�&ni�~I�5b��j�M�`����}���鞞^77�@-���Z��XN�u�Sƀ޵�=}�1�<��'�X��ĳ�~�D�1�-Z*C�$I^8��UT�^Z�?�eb�|�%�?}�4koi(h�K�pZ��ucHYz&�Z�ɮ�h
�"d[��=����'�@p��-���VA����ժ�����IC�����:6�g� ����v�*�i͚O�OK/�?@�Ȍ6s�jR�念\cֈ�si>�,m��ѓ�)5�����Y������Eù�=����{k��a�j(t�	���R��j��K6HWٴhZ�����9����}
�G>M�=Q�ӳ�q���y<�⡱�Yx��EFOq�N��	��n<�:��r��K>�Q=uܲ�(�Nr��I# �rD��R�i%���կ���UC��Eg<�
��@��H��"��Va�J���}᭐ІM�����<�&��2�H�ť-��n'��s��嗇�t��-�H�\:�1�(\7����ď�V�^|�%ZǑvN`�ʥ}��Y��Jwu`$�M��GH[�/5[hu�ʹ5��0P��m�� 0��t���e�ǐS휜�˸)\]��`˸�]Q�������/��h��i<b�'��vdAG���+��h�í���q���e�%��l^I?��H��r#N�+�`�w�W�TJ�T(�t ox�S|(��*���H	G�f<�蛉�ͣ@�6U�S�#��!�tX�q�B��S{E��mu�l��˧�&d��?V\���՜�_)�S>vr4=�'3���H�MԆ������j������z�M~��OSx�jy�֣�G��m��0��cy�XB��Ǹ^,>�l��I���E:y��rǙw�<����s��%�o�s<���ETiD^R�o/��Z��WF�7�	<�t{-2@��:�V��Ώ�5�["��a���6M�]����W;����}�rC��=��<���B����T�~뾢��+Ktg����³h�9����+$��\��!�2�S�w"�D��u�m�=�Ğ]��V�ĵ���cl�6t\2��A&+���< �[��f����6�@�����q3��q���!��߇��τ�.
B,���NdJx5�>�����s�9�i��C���v��l�0��3�۲rV�����!�l<x���隥�쐊6���=I�6��~Z�#�
OZ�'��2C˹���W$+���z:.ӮJ��!�>�W��𦸵ȟ��]�7;�r3v�9�f�ˬH��\�P�^��䰾�#�;�w��B���&n�������i=�q�V�}��"$Y͑O3�M��c;2<��\.�Q�3@J޻�:��m�.�:Bg���E��b����n�'���)�Ma}�Y_z+��:gW�~O	�����ًɿt� A�7ɘ͸:GH�L0�8�,�4���"�tzYr���V,\n���+ �D� -^J�4-�:�ݯj�*/̥��3��a��L���c8Mw�"�0����n0*��/�=3[��`����m�Q�@RL�����5���w�`jøn� ˓���t����t�뷘_Ѿ����ʼ�r��{���j+�٠��m�0g�2��|�w|xhP���FS��>�ҵ���i�["K yzP�&��q�=�����G?��yK�Y���)n����0C8����J��/{�� 'Ɍ:-\Y8�O ���N�B�
���sz����c3-�F���Ua\;oh���YeUO�f{�	&�O��ٶ��"��Sސ�ָ�{&�x�Ǜ�׽������9:-x&�;�V�k� ӓ���4QS4�rP�$�*ll(��IK��]?�R���ȓ��*�W�G=+�Wl6P]n[zl��J̔C]�=���*X{r��FjLaC�<�K��v�0�j�|4��|�K�����>�����m����J~�Di��f�!�P�q��3��5�T�
>��bJ
����W=�	��=q�8�7���6��K`��U�m�T�0�B��x�m���>V���@�CZ��2���f��+�)\˯n���|�f�_s����̳����@h`.�k�X����~j�/Q�5��&��c�������A?�4���e�|\���M߱�0�vN���2d$K\2#Xks}Jz�n(�$���d=p#=�I�i~.�yb#��v�w4��{`�3�tI"N*˒*5&��U�9��h�n��_�0	���� Pzu\�lWn/h�-�,����14�R^u�����q�h4��6mR{6�/ņa
�qkc���ר�r�(��y ��-%1˯4'];�4S��wJ���2K�l��@P���Az4f���H�)�  ��c��UP�c�%�V|fy�j��nn�^,n��bR����u�ྼ�*N�}4dEyU�_7�.��{O]�>݃�8��*>��Mw��?�J��kb�{�t9����� 5e�(i?(��:ވ���TmuB��Ƅ�����YՊ�6�_��tF��̯c��R,Ym9���{��O 6����t�	y\�ԧ!n���	��8�4����(�NA�\���y13�S"\�Rk�b�����Xu�:�e��k���Mײ+BQx�<�4Ģ����z��Ew>��?�����)�F��
Q��k��e\��$��d����F�ǢK�����v߳_�i�c�~o�.f�U�œ�Nf.����_���P
�%��v�<�v����4+&��V�v珙��̳츝��E)��@����r�c�V�*�7�p9�~���^�w��;x��6jH>��{���m�R.H�+����V`w &��2���7�u�o����1}�u/8K�4���۩�z�B���ӂ������6Q�<��u�#�M<(~,`�C1 �����T�c(�C|��2Tx�*�$~�:���؈|�R�~����^�{P�y �W�W���8OK���Z��v~9����^=�k�qmJ��,�_�
x�+@��X�zpSN�h�����N���v%�~�S_Z����l[07����	�ҹ�3��0�@�Х�zG���ZG^�s8H��s %�����G�Cr&�V�&-��9uvQ���.�w���e� ���5��-.٠u�+�)yx
��NC���c��FD�Ip����@4�����[�:\�-��� j������,S�c���"��Q��THK��{�2�[,ݾ6$��e�Oy�*�8>��5�a���V��S0��8q<��L<���"�3���Ȏ�=�����a;��ɷl0�@�!��1W=�nB�|�����y$�o�e�[�*��9
�ۓ���v�����D\��1A�(T���_C8��ǣnk�Q�����z�6 �n��%����c���E �f��o��[)�;�<ƠX�%�j�}�x��
�mWc��w����-��S[��Ϙp�H�.Xe��3�@�.��F�����HCc���*�n�Z�t�%.��᭣�Zya��ae��q�5]�$l�F��&��⨛�I,�E-��\�cbX����o���S���?�QN���Ժ�ks�FHRl�j���Y��a���+��<�z`�-�3j�ghy_��Q>+�PgQ��vI_��b�G�u>:�����W�9S'}��L;���u~��,t&:�Czh��A��?����龜����옸��EM��>P�U����	���%��6x�uN�c;@=�
F[��1��l����2��m,�����Zz��ޞ_n��J������߂���	j���NC�b:%3>��nH'<�z��_a�����n�J�������3��z�����NJ������v���a�V��!��(����N.�ܧR_@����ur�]K�Հ�N,��N/�i����C#�ZgL($)9RWH�le���z������'�����J�B���z�ݍ1p�N�c�����Y}ݣ���K+�xj-Q���� �)`3d^���LD���^{Ę�
Ÿ6�!~m������Pl����D��聕8$���<ӳ뒝�P�����C� -wo�p��� 1P��waq@PS��ߺǪ�-Z�e�{���:��=��ۀև���+\�1 R;i ���"6������"�/�!�WAB��؂û�����pk��<+��x����h�mI�+a_�6KG���͓����]m�bd��҃wL�4�
P�v�ߎ�M\?I۬�ߥ�����)��K�k&^c�om��$8���x��L���5$.P٬	�0����H���	_��/f3ҼU�+���	��	��ՖM��񣅹x.������Ā˩<Q�7�6�k�,��-m*������C�!Է�~�0��AsKDJ����!���֝�)��_�P?��_�����g7FH����}m�2�)�I,w���v��݇+^�˱C��9Zq^1zQ,-����)B�>��U����"D3�x��C����_�������m�S��K�������h�aQ���ߝ.�����s`wu��aٔI^V��r@��P�{hDw��ni��7C%��Vϵ7���f\z��� #}���&�*h�k%�o���kR�\��i�
c�i��)��Wzw>��2�AuXg����i)�B3�(���~��a���Dǳs�]��"�跎U<p$g��˃!��Ѿܳ�G�.�=Ui��@|�̜>i�tB�s���5J��l
_}���rE�&�Zh��'��	'o�E�I#C�;��;$��|wY��V�?��c�8=���My-ˋ��Ňb��r(�������
�2��2�����r����wg"�d��D�Z�<x^�W5����i�^�'�~��]�ܯ�a�-4gVn�k䪧)���4��[�4���
�m}:��O+��6N I�꒸zǑ����A:� ӕ���A�]��#{5��AU��������mA0q�ˑ"�Db[7f������L���gMĨ6� ��	>�&����	d�'j�G�P�Y�uŞ9�X0���LjP��O�`F�#-��9���ZOB��]��qχQW�a�h�>%�w�x����0�?]��B��NB׳2�jeo|fWج��$m�zL8�8���傹�]��'�ý��|���{��~	�3��9q�sH^��1D)�	�b_V/�5��{�L/�B��O���u�����	�a��D|�ޱǉ�[UW����.=3������YY�֨��D
r7��߁�__a%cup�(�?Q���v����%�5�v�[5�VR�%���w���]�����������g�Z��r������B����Qz'�g�gәF����&k������[��+������+�NV8�%�+8;R��h�>�ޢ=m�KK����Jĸ��Z�.BJ%��U�vj/��^�Ul���s8G����ܦ3�c��@�^/:-\��k5�{.��C��rʩ�֬�/���ؓ�������(��{�����L#�WLe��o��#��3�Qc��Ӕ�$|3����Ck�ˏ�z��woGu/�{�͉@XB���חS��d�lr{u2�0.݀� ����#�=e���6�u��t�?��^r��ׅ.hOJ*��v�Q�a��!������\���Z���zr�=C�ϋ�8��J���L��$mK�	�M��u�Kq�
���r��?�/١+��V5��BOW!����u�!��=�j	"lҁ���`�/����)���Wf+�j}4��(,)怤zQ�;�a��� 6a��7R�"7�����z]`��gϦڥ2��#�K2��R8�,Hb�b~ 8�,��2k�+�ئ�ү����x}˒�����j���oy�h�j��\z�i���*�����+��I�<Qh�l�n,�q"�)�h�y�b+�~-v)X�v��(+&���U�މ$,z��˖�rM3gֲw�I/�
��NN����n��-%h]jah��L�.�rl�5�@\[��B�0���޳�?YvӘ3@��ϛ�1�=^c�w��O�~��Z6��H��	�]5�T ^�J�b9��o�0p��/{�!��R���Æ�:��9�����r%�h�_�2!C����.��aNw�o�8|P�,Q�-�W�����`�e��OU<��<zE �.����1�D��N������� N �:K�d-J���s�X�ǩY�R���<7�>>`~jݬ �;<C����߳��������@V�Cw�D�� �i�ɉuA���>�_pY����n0ѱ��dK���zg��|�G�gg�%������瀢:����C�h46��wPa�sML���.C��oQy�ޤ�lmBF�X��o�+��D���y���G�2Y |�k����w����"/8���`#z�1��E:?�.��]v-���ߔ���s��v���w4�<�eWg�?�OG����M�*D��	�	�X��n<uL�E7�eJ�0���L��̣E��]!7bQ{��D�@��k��)����u� ^!�J ��{`e�&�צjPHƄ`�� ���ek�Tr"c�Z:Y9p�������ο�D�|	BC���[mת�%�Q<l�.1�	���	��=jZ����� !����������p%V��Ȃ{2L�W� ����w @�e�0�Ճ'�  !����Hl� }%��V-Μ�K�dM��r�jxj]�Y��!�� ��a�y��}���<���{G�8�gN�����㗘��mA�oN���W�R>^V���c��Nʊ�v�Ʃ�W�� [��p�o[�9Xԝ�4d�$ߗ2;���K?�#U"?��É�h�& �!�3yh�t��'Jb�3�����r�3�]��� ƽW	?W���F�/���Dw���y�f����7�R��W�X�����V�i˦p��4�)5Z_\��O;`�n?��M8�2�#C��j�|'2�$�L�$A��/�\���hMkܛKe����9�>w���t:���PQ���Ć�9t�5�c��8��x4D��]���>Ϛ�SnepK�n� c�T2q�&RA�au����;㟚�wm�#냸��5�Q'D��/L����h�����G��c���j��<H^�����ۛ�D�,ub���v#PE�\�IN�� �C�?ﲨ�M��2���������Mg�z�j�'Qv�X�C�$��b2f�r�voX�P�q�x #:Y>����7*Ȝ�k��9�Z(g�k�,*��n�I�ټ�cT%+�8��$SߖbX{*�'n޽�p�, O��������W�h��I
5��cH�	�leo�Ff�>�����'� �M���e~P��G�2��1�I6���N���]6.5�s�Er���W�I�t�B�+�?�}�N�'�	R�<���go���;A���q&N��t�p�	.ţKHjhV6����S5��6Q6{=4� p.O��U�H�����J�>ݡ+���/�p�W��8_�žl������`�'�f���ζ�)�u]��A@]��Y� .+@�����q�Չˊ8F�V(��$��
P��=?�&��N�|��
=����ey��*��3��|��mrl�<ɝ�����9���N��J?����X�H�m�L�̬��l�/�)ܖ�nTÑ��+���ly��ﶤ��o4����oe}s��]O�9�ԧ��M��L���A�{jм87`v�U;qY�V�S��B��wN�
p�2��]-oD5}eUߺ�[��~W~H+�:A�i.����N�b5˺��Vf� ��X5�+?�U~�x�4Nw��[��Åμ���n^�I��0��-��^Sצ��?5�R���9@HH���2ܠ/:����K�=u߲�����ŰgZm�d؞��@Q\�@���
�v�I��[(F���@L�AC����z�J&�z�#-�f�<�U$���C���u]�������M|<O�@jLH��J�'��>S������U�$��N�?K�L��Y?�-�:x�<�^�` ���sb�H86$�`�=o�D��D,�����=t��S��[�3�x{1I�s^�.����Q��=QI�q���0=Π2O~ȃ�v;[2Yҳ�b׎ȀF�?'x&�EH:�<j<�:�u����0�8�L�G�ηؘ0V�=M��<�c�5^�C~S�G���v�_���+Z�����h�p�Ŗxg4\�r��~4%G؛�g��{���ng����m�I����i	h=�T��m�=ώCR�5�3q��!On��v衤l���]����W"�WC�E ̾��Z�=:������g��V�m��x��]��!���M��"�z$�!�qג�3u-����}�kC�va�=V�泽�Ь�,�����S/>�9zj��\��nGTd��4�?^������	�;�=�nri�ə��I㧐�S�Bu��(��[�?[WW0"��2A����I`��sһ'��H� ��svt=*[�W�V�)��(�[i���@E������~U�H�Ʀ���4���Q	Zƃ_�2(uّ�}����Zٶ�ƇP,�*���}-�-H��g�6��oL��DG;�W y3z]}X�Q�Au@��+[�E��Պ�'����.|`\F�ߧ<���gHI,]`�_5�&5T*	y.�`�@�pk�QC`�'���g��%`��	���y��*��Q5�Ŭ�O��"��\5�}�O�LZ���/��R�<Ǚ�����Y���&�����3S���QK�R.e#�u�ǽ��Dq���T,x�s���q11����f�]�K��Z4���}$��ɋdPd�	�}�`}�b-K�tW�o�w����H ��ߌw�֨`�(�9k�R�^N�����F�KRj�T�>�L���rn��F�g�q���ގD�O=j�TZ~3�3�="/����N�x5��������jj�@��("�T�"�;bA�Ҥ�*���(���B�J tE��4�I �5@���;��{o�;��u֚kι��guA���:
���[9ILay����Y�e��~�x���� �݀�B��lxE��
;\�tV0��|d����JF;,N#���#�k���?I<�\�72�5�+,�UX����lW�LKvҩ���*�eC��g���Tf ��Z���|����5�z����l8\Y$o��D��C7:��P����V�b�d.}�,�	/�啿�t8�����3` kTR��|>8�տ5��ok���~^@*-����{��P�n�km�}��*TM���>m��>��r�B����V��E]�\Q�����E@DX�
@ح�����U��^�sBo���� ��Ҥ�b��[F�L���0Li�9}�T�#�,Y�0��T*1�ߪ���S*����7G��Qe��*<�*�b8�� �7�4n+��dOU��	�QȾ�K��#�����초�J¢��t�����#3�K�b�j"R*/d�����<�_y{��%\K�`.&�*� �4c/VUA��B��U%����;�f�=g��1��fթ�ˠRl�␆�V�VG���v�� Iqm�r���y���W!"c�3��6����}V5����H�E��&�bbc��~�{���Mfz��3S2��qo�Y��rNf3Kvro�	�����em�!,;����f&н�>A���aM����(���}%ܨK^�hL8��'r�������i��
�m*��#�ި�xs
J>�b��џC�@�(`���*0C$���M�c�N��d�72櫵�o�/�ha�d$�������R��VX�*˜a�S�m1���i�%r�aV:����]y�f��op%��P����"�<P�͸�?P�>����kl��[7�&f�O����4c�����O�,r��wk�%.��$�eB�ŀ�'����O���7�{,��t7��fÝ�����Oob�|%p7��%���=[5�~��1&�i������A�?�X��!_+�'���Co��6̖ȷ6���o�B���^�6
��>�_��48L�`]u6j�4����>91M�D�I��M<�It�w]0k�j9rf�D��v*¥�DSlM��T9�E�}�I��(OY	�n�J�N5����q�7�'N%����0�Z���:�9r���+b�3x�D.��<����G��:7=t{���.ѹ��	��,���h��YҺ��,��&l���J�����r0��̮�N���"�>���Y6�x���i�ƙPAl���g�jA~�ĄK(�z5��'S,~a�ɢ��/[?Sizf"���ֺ\�<U�:�I<�cP��6:"����+�x^7�[�TafM���V��)����g��R6��#v2;�m1f�E����9������2�r�Na���?N_?�q�����݀V`�o�E�W�943�(���s�ns�Z��z>FB#/�efg�7���A(���Pb�X��.���K�÷�N�??H�"�����9�k����+Z�������ŘE:ঌ�y���G�$ۤ�ڋ]<Y�c���T�4��vP#��!�Ib{��Q۱�	�7��u7x�-u_i���q��9�4N���$`�E�ǟ��wZ�M�L�� ��1� #Py���b�М��Li�z���у�-j������[���5d[탵���ӥ5 ���w 3:�%?s��O��C�x�j�E����'~"�^Ti��H��7]<5����Җm'}m�=��N�,HU�2��*`o�Ԧ��:��Ur��hgw}��͍�!'F4qrnI2`��,���{CS,+W1!b�8��(*�	 �r�����6�x,c)sz�Q����>�,8X����f����Rk <�]po�����u;V�X?��S;���߯��� -t�g�?D�#pyIm*�14�W=�%����:��B�
�fꧢ�B�WO~��d�_1��:�CDe�$X�F(*�c	�)ڃ�,A�]�����RR^�6��䈟BO.�t�=)���'��H�Dj�eK}Ǧ!}\�YX�qq�K��̢:��30����x�
�䇻)/��$[o%��YV�w96�g����ES�os&~a���2�.9&�f���u��I����o���/�E���o��;�n0��D]�v��"G�'�ceKp����g� �\��Ԭ��}O�$����R�ud�Bo��m'��@Z��p>m�tI��:�/k\@����~����,�`��i��l�%�q&ދ�87黊>�)�5��G�!i�S��1h%��Ƴ�/�� ��dY��v�|�d7;\Us��l�����f%F>Ӕ1{	1���9�C]��mh��BqӲ�����7ַ�������(��@B��U�|���{�ؠ"뫺�TBj������WS#���3��Df���E'���O�f�N
1t�K�RG���G�t��6�O�V�L�o" q��q���0�Woѭ�{�D��k
W��Ơ��?RY��*�
;����>M�e��s�-�lc���s�1V��3~�̫��o�����r�"���N�i��q�����NoB�P+�Qof.�
`"Zش�?�w]X�eE���`D`��r)`������j��)V�/+���>t�>Qi��L���P���J4������)������12�[Z{n�	�B����;�K��"�<kۺ���\o	�f���� ��4=���q����o�=��<����j�S��	��}���̡M;��q�����]ٖX��Jgk��05I`ZykH�[�=��������ɭW��g�vb�	=K=�aq#����zY��G+�sù�1C���O#��t^b��j�	�����rBw��5��/�}:�X�Wl��E����J��\��Y��F4��Z�'V\%���y�J�L��W$�-���y����ܝL/2/g�5[�;���¥f;g�43�'�Y�̵�����ɎN�#�jR-|�-)o]��!�E�'��D��D�0���1��UҫR�XD�}e��68�����Hm�O �}��o�~{�L��l��✢�����-��i�T���cei)���[���?�1�{�4v���ӫ��Z�|� 8���絻�mC��|}f����g/D7{��H��۟O^^��E|Oemym��D�A&�A�oy}-N]�?͛OZ��jZ�n޺EF�!�|�9�X_�~Z]���MzEq�}~ƭr�Lb���㇯����=��H��UI�a�8�S��p�E��e5�g,YǮ�Ȧu� ���~�?��{'d�f]�ik�%����Y	��W���ZՉ(�{��0OCYD��8 �y��Y��9n]��L�
3��+�6�)���	a�m����>y>^`��qKͳ�q���`��䐩���<��Dh���;��n�e�ن�òY}7Eo��e�Y��VG�|=b<��:��g �0t�"��E��E��F�X�8�f�~�d/FN��4au��.ax���}�+W1�vO�@ȵ����q�h�4��;�o��锪H�0�2%ɒ��$4�	�y�fG\:7�U�����r6����t�i���w�*~�H	�V�/r ��w�p������P�d�ݾ���p������r�O��dפ��uӖߊ�O�������5e��fB�p��	���"�m"�F�y��*�/m<��fI*0"�Ts�寑��B�`�1�P�KXy�}���P�0�O#E0�/�ˡ.��g� �q�P�'�9�+����/��侱q��5�.���%
�1�� cQ�^�����+m�����!!Bh���Vl��6ǁ�,w�����Ŭ�,�m�nc�-0i�3|bZ.��n�&^S�'=������2*�bF�ҙ�S��X'�Y��[�,��h�f�cf����Yz�%��ys[�W��B2�6�0*��-�_<�8e�̢!D�M� Mq�H�i&�d�Z���]�pF�O�E�
�:��EN�����%ͩ^�Q� ���N��;};�U�D@�2���9�;�8%ɼ>i�.����*v��X+l�r�-7^n���1�V��֯d%J�59��WN�j$N	��+%R��oz�%6b�_�O����o(��L��^oKB��[������&@�o��T�֒P��%���B0���d|w
��
�Sl��$�������};t�f�jS֨b?�A�c�ڲJvV�D?�F	Ȕ�<H��m��&=�]~�v�ݽ ?�Ǵ������Ȇu��<ƺLB;��>�Q��I�S࿸rҩ��e2�=��B�0![#�͘/���WY1���r�C�[iD�$��Q?�B�ڹ�j�P>d�Џm���B�O+y�w%�.���K��馮��$s�G	�l�{��� g׾�V�^�i��d/5g��|T�w~�b��W7S�� ��	7���c�}�2����/�X�G系t��1;x'7�
r=�N���U}�����G��l��#��uC#7r��㱳�U�6:��s��|�2��ou넺 |��[��-W-�)�&�\�N	~ba�/"V(T�jQ)r_�*�s�T�QXE�J�v�DdJ�E9oy&��)�� �����l��H!1#M�P��tr>Њ�295�T2���ϯ��r\�����(���u�o���ټRhrT�Ќ������ �YF���"5L�ɵi�1�uH2tB���aL4��5����tk
'�q��w n�%���?��}�t��˶y��8I�H���_��ۼcip���~d�li�M�����'' �CD#)%{��
��>*?O�	H0��v;�Te1L"È�.ek�P�y��_j�Pv�`]ϒ���WM1�?\	�ufgb �`J臇d��q���vqP�K�P�hOF综�!}�K�(�m,�M��k�Mgڨ|��m�(i���Ϸ����R_����j����	޾�,�^J}�������5���U�:�+�M�k��A�5��~����@j6rß�L$�16�o��E˾���k�	Q]���E3l��닐�N�Sm�O���U?Y=1�-��Kt�V��c�4KX}�护��J1��sPg7�j����n�g�1?��N<����ֶiM��}0&1�q�6(~Jd����ط����9��)��8Ó�g8n\�N�#3�nqa��[K�V��vXhA��%��FK'u�ej_�
گ"k��+@�-ق]0��;�.��*NLB���SR�T#�WÃ<8�n���/��_�5]t���;�4
9�r���<�fV�#�����aH���ǔv��i�}ָ��0nM��U^�rVf�"DT��ĂqpV�_z��^��%���ʕ���ɽ;��	'��1ϗ�6@��F����ń>���GnѤ�p�!:\�d7��rT�/���ҤϨֵ�z��ࢄ#�دԓa�j�[�yfgW�xV�|N7��� ���h�a�a�$4)i<����}gj>��Z�&�՜Se?A�h!}X}�=�0��Y��(,.V%ǒ��R�[^�՛7p��%��r�������,���w�e?�ce�e��&�p��j�̰g�y�#vW�u"3�X�/r�pc�z}������Svsd c����U�ԫ����9_%Ϛ��|��RkQ�����( �72��Ez�|�_U���������F�M�}8��Ԍ��8�'���}mb�?4k���	hf��3ϣ���b�
uI���x�G���=��.�d����uAw�ȑ	n2��������O�r��0�oago��Z�u�*޼�K=�G�@���k�a1'}�'�<��E�w�z"`m�ˀp�V��Dq�ʝK��3��b*Y��)����,~*�o �O���In�f9�e��#䈓zݚ�~fw2E��x<��������g��_ݯ�F���U/+�RQ~S��hB�F2�W�K�#r�������S <�Ub�$d���l�Ve;��a��+���M��l�;�｡O�8�����������������ϧ;7�He��=gdv������C[�DDv1k_P��
d`�W0�����$8<,H���i��[{��b�M�k��j��4c�u��2�ך�̐7��?^Hª��<�w�,���Cf׏����(�m�\Č튂L~����\L�W��X�@G��hx�[|3(Y_����z�ȌNd�*��ܐ��.S�4R�8�q�}��ܸ���3�,w�T��?����� %g�%6����X/�v����%&7����K�g|��EN9D�H��i���9
�N����~+��
�0��J�Ӟ+�+���.i���NG§SQu#ē���2ua[Ȳ��yʐa%\���xiI`�1~P4:���̓J�F��Ϛׅ�٫M�m�n:��/N>�>ўJ�?a�t�؆�Ψ(@}�	�a�i���}d��;�U��O<�V���9W��䶊��LJ�i�1je��˓G��QE�ޱ"c|w��W����b���>"]h=��q�\��j����?�5k�Y�=>�ɶܳ8�����S��e����w�2����X�S*2��_��+4E_���w �p�\�t*��GP�V`<�и�$D
�p�i/�&��a$��BP�K���W۳U��ޓ䈚Q[��9�߮�L���f���rB�ēq��<��8[�MG����@�!r�W���pV}dn����D�yS���s�T,�d���N�§ᨀ>�O���ra�|����11�e��=��k��*˱�{2�`qC�vgP�� ��sw���X�ɾe�B
�nX���b��nv�¬}����[1K����>g�[Q�쇯y�z%�#��.�?bb���P��C��E~���br��cE��di��*ٛ�Ќ�i Z=7WY��]Ɲ��j�0��5 M�Jq�t.)%�H�;O��y9>Vh	5[v�U3J�b!\Mމ8k/6��ء[1��%�B��ֶ|x��8�\_�T���mx�����|Cv�D�c.\Y�H�^īkW�2��T�sI�tr�O&Ja2ή���7���鏉��y��$/׌��{�s�}\�W��-p�	��v?W�W���Ͱ_�j0�+5{X;��X�UG��� ��-p"%B%]����-̋w|�2�`��<j�pF�+�֕s_����Ņ ���ľ�D?�؀X����y�2�*w4y��`S���!�fߨ��bb��	�Թ��݁j&��yj�2TZ�s>�E%̨��Փn-ċa����*�B�=��=��P\�1�orP�è�m!�9A�	ΰY .���㯉�X�*:�̛�����Q�DE����/�[��-�WȓW�$��c)@ �a�T�Rp+�CLˎa�O0o^\T)#����CF��X���+E5G�����SS�I&*���Cw��;W #�i¥��6!\0ܹZ�N���$���Ơ��*�|�3���5�R�r��t�@(���}��ɠ?������}Bش��FE *N��m�5ZF���Ci�6�*���� �M�P�O6�-W%W2�"fb�\u�| ��;w�u��g�2�]��Y�
P�T�Ҙ�֒����n��jb넴[~�ޞ�x<J7�T{�RHq7
C�y<D<���"������ç�N�����أl�D��QLB����%ꂪ���n�0�6�j��_l*ԇ0�*��e��I=����M,V�:����U�\8Q��kL��_�����F^��{����7�L�p��b�q�$o_E�"���y�Z��E��x�yb#7_��mn�W�]�����9���b��~���,п=�L]2ޱ�����%��',���J�V�F�r�%1L5|C��g�,�v��o��G��bCjfJ�x��}n�tkH�Z�p��u<e"�#�E_SɭA�ܓ։�N)���,pz�;�h���]�(�?������0�����B�te�
1���s�豓��"�*�z@֖|UTҵL�0_��)���əqI#��_P�S��N[��ҩ�fG���|9�^M�����P2g��V�e�tw�dn�I�2��M��9��/Sw��G<�>�X�"|��7���wVleW��cx�*f���r¶yf��$��=���;5��:�4����A������_��%2/Y�I!/k���g/4���?i9�8���jSA��<��NxAU�����\v���o|)�j���`/^��e�k���_�;|;ґ�h�0ߪ
���z��^�y~��� �J0xqQ�W�380���B��@��<R�2�8N���2R
5 0��uab��zz�5S�8Z�I5P����CnUǈ`��b�]<��@~�Z�ŷ[z��p�N���˾�$�O�E�/��|�?���I��ɹ�P�7�A^Mp��y��9��d�P6��4�9���.��įx���ǻ]C�Q�q[{��!���IR��)�P��K�x~�%�oę[,c�����T3hWa}�;����#�Igڹl|���H�ߏ�ɵ�
y���Ќх{�ฌ��F��kB+3l���>�#J��~��<�j�8BhA6<mKHˣr����S��	��Ҭ[�s�p�HB��iN�@�3~ь^h���k�+�l�[ڡ?y�q��EK%��_a�a@	�`C)�}4�P�W@sP6�@���.����0!�4�ui�@�r��m�j?���>oaaЭ���
P�K��H�]�*����$Nb<��ל;���S)fM;�l�YDCʢEޚ�F�y��T3{O�|5
���]�x�Y���e�奇t��;#q0yO4W� �t�ldkO@����+g�����ch���xa���� ���7;J�sl�x���_�m�
�Ҭ�d�:��)7�a\bO��F�2�w�:yX��H���r�������$�U�u��Do���d���ñؽ�z�F��64���6^G%U��6I��0�~���t$~��#m�݌�*�3�0ް�B!G���~��z���%.`5n9S����lQ[Z�F.�{��^�{#G�/t�c��҃o@���|-�ݚ��l" ��O�5L� ���0�QS�HQ�I�p��Ϫ�خ�Fp!�D!ZNŰ����{cR�=�]cvv�w�n{��);>��<V�3f��
h��w�}��s;�;��6&�2�\�J^Q�Avr�\m�y��{�N��g[?l��ʎ�x�:�7�_���ۥ�Ќq�k��K�Ϯ�?|���ɷ`��#l��ù��"��n[�T��'�`xy�r���,������W���ssv?:g��E�A+���I��������Z������r�Xw��f�1.I�؄Hμ�u����p4Ai!Yi!�1��]���Z��������u�������9� ���1s�ʿ��-rv��S���*껅����%�3ܺf����d������w�n��ùӥ�6v����иפ��v(+WJ���8�-x��B�6�RG�X���Ќ=4&Ո�pv�]�򗻊����R0���.U��01s�XG�������py��/A �t�.�k0=���5MI:H��0�~i�Њ���y��x/n6�ܰ\���W/˝aͿ��x�g��Wz���% ����z�)�@�ӿmg5�j$�٦� W����G�Pʚ<�P���.˲:nq7AX5c�,��ks�	32J��m�Dp|���[reEo|~�h����Ѹ��C��0��{@r�3�us�ސ"�6���G��R�k��C�ΰ�'>�j῏���6��Mx�v����ȟ!�1��@K����RHЦN��]�/7ļЅ�k�2�bgWU^���ԡ�o�+��t|�0�!���[@U��d��I�X�[�s���A�7ee��݈�9�gOU<��;����Ƃ����c��[��2��x-���K�J�zt���e���m dF�8v�O�TR6�đ:��;�1�ϔU/7�B�o�9X0�E������n��lL��B�(-{2�c���%��@�W��10Ψ���^kvy�q�E�.|���ؤoRh�Y�e)ww1Ŕ�˜�S�J�f�kRY�@^��)�MSZ����H�+���$����:*���d1�R�Do��q,��kE�����@I�o��D:����!: w4У�� �E3G�ۮ�1�.e��Kh��`���a��S��\�4�8T��;��<����<����>��T��ާI3X��Q{Q�xT�#}#��\�!��w�C��/y���Y�E�u�U~ä����n�6��ֹW{==�c��pBQ0���1xo�+g����P��L�����}�+�^�.��taey}�;����-�7^�{ߌ$�Vi`0�z�ˇ���[H�m�7�>�I�D�I��ҷ��%r�6-�w+����!f
��2���1<+������e�Y��� �][����K�Wjb�� �Z�Z6x�9����/����2��K��6mM����Fș{<E��̂���K����vЩª��B�.T���TU�m�o����@�s��t9{l�EJH}�݇���n�&f#PP^��F�����ݓ���m~ ױ�@X-?�8u�<j:h�7ӡ���=#1!ִ������r���ϰ �[�ʩ���L��e��KP�E��:����uvЫtb��q���:��'�hYL�!-�X�({Z� /��y8S)�����8jVwB١v/��j5����b�(��tD~	��e\�z����B����jYF����j9����<����#�!%d�İ���+�r�:V���ހlf3
F̥�j����� #��@{�9����lj�fŒRf9�Z����q�!��!��6!]�wb@�vA��4��Q�@�G�!��z�@�g�P(��gK�v"�<V�������˅�̍���R7_��X�;>��L�D�
*�S������.	p9o�+V5��{�&Y�@�|�.��V�`-��#����B��0x��AH0w[I���?��%/,t߫��>�o��Jf���,�Y��	��!�gH�d1{@%j ~�'� ��N=J��,��]}���Q�hzupo��mGJ�֚6.���e!J�&5YS�����4�,c�tSK�Z��^m��%Ԍ:�-c&���|���N	�S�O�~���Wv�^�(R���y�3���l`���y.wNy��ϥ��*��s�G��I+��>2��ܝ���},�?���_oX_P�Sq��(/���	���J;�i22�h.���FMR�]&���*U�T�T�J�퀴-W��W�����e|m�̤7t���mE6(�SRd+lb�3NRk�\E�j/V`4}���yulp�|���WA�mK�;k)�����"&� �l��,�f�t����� ^�s�PDp�D	��T`hM�&mp���n�F��#����!s�j%%�����Eڪ1��%���ֆT#����Ȇ>�X.�S,6�lI�q<�o�2Xz�(���
�g�`���<�
��/5�[y�B�8o9c�w�˝�\�\"�;�Kr�-�ՙ+5d�ac���{�U`���jþ)g��x���J�&�<Pe��8�Uցݿ�?�G���,�/��^��J�O��n:�/r�]jd!��_���9��
�H���W[�!+��E�/�g:΄������C��m?���ؗ�ˌ�l�W�6�j�q5|�����Zu���P�هe&�j���dk�K�O9f�W�������!KX�J��4��{9&w~�,��*����H�[Xz�����)��@ޗ��-��65E���L�ӛi8c�iA�~@�����;jl��|f%_t	�+8�����w��s�WF ��kw0�.�Y�߻1!�m6��7fS�Ў"�>����:E�[\���|��-ēf�f6R�R}���ͷ�F�QE��A|�Y"w��O-pN>�gHm�;��40��x�Ӆ�G6'���	٭�c���6G�fv#ͮ,�_�Ϻ�M���0����/� h�ΙJU7�,���Ak�������<�Ut!u�P5�v|M���w�hϽ�ߓ�E�܀ ���{�>����'�]��G;鬲�]_)*�E\;�5��9|@�=sѰ�m<�ou���;�j��#���Z�>�]��2��`:z�ײ�W�����:�d��T�n 8�EE^F��^�j��� ' �p���|�3����>z���?�g�{vr��g�����}$Zη�N��~��oy�}�-{��QC�_�;Ě�Bhso	�Kz򊘦������]2`Z�g��Ϊ�:����ɐ断,��;���yoDZN�h��>�X��ԐHYz)�zBҸ�0��m1�.Tŵ�O}D�dK�������^4��NC��X�1��[4��ˀ�y��m�憌޺xG�?���*�l�?PCC& �i�Q�c��栙Z����*��V�x��%T^�hs���b��پ������,�׀*ѵ���|5 z�� Mz���d�u�Q�,�r��b�ю�
�����i2ސ~n��d�F��_��Fq�=4�U%�xAUf&�#�'��TV�[y[��ˋ_`宜!]�F�?گ�W��j��Id�&Ot��}��ꂈjM�<ŖGC[@����K �A@?v��r�bYh��Ddo�m�ktOet�m+W'j��$y��uSh[~���_���9����𰢱���U�^D�8�T�MbdJuY͍��eK@\\p�anN��x"�y�HJ�Q���5�SS���Z�?�ɗ��^y�<����29���!��Aࢋ�M��C�J�3��)"��>�8���*j��oI.�q�uβMs�3�F ��3��[OZ�5	5b�Wɾ12�
CC{ �a�bK�{a"yo3���/����?[��o�[���c<E�~��)�QΡ}��w��>2��@���0�+����s��e"
)������8N��FC�,,��]:~�l(Y|�����/|5Nf��Z��Î<��gR����z[e�k��0I�Ղ��X�بʇ�, +�q2��������R��kB9������Ϊ\b���Dʺh���E�A�Ke�{'אw�Y�Wߝ������׋��cs�����22uaZ���ں�З~	���v�5|�T#~�M�+���F�M��^����[[����A�f�����֝Ҙ�¹�G��֝���
���0ghxJbڏ"�n�u
�� g�eV��&>}a☛�k=(B��z���#}�r��p]�9����nm��d��A��q��V�<=B0���	mA�����b���T���XhŦ����P�Q��g���d;�e�+tm]M㠑'V�I��V�g�.R@$�˯	�$���V��,�/�d/,���p���ھͷ^-����=$��Ok���XH�H��O֓X0'Sm�֟|��O�Ξ�81�
�.�Ӟ>i(F-�V,Nn����?�c�"�byN(6���2�s`�v��:`�K���Fuӟe�m�A묚E�a��X@GJ�����B��e�E7,��t�T�Ƙ��>�?��d��W�l腫�����=�z�����yEt!�o�GJ���l 	2&~M��c� c0ѩsk9�E��J��M�o���U'ځ��П��J5	�c]C4������
�^�ϩ�����~���v�/�d�4qn�E��O�X�+~E�z	0�3ߋ1l<�7�LI"�:��S+ڟ�!��4��jӽR=Y|�Ӳ,��/�^�o���H�-k�~�y��a�����zZ6�?;��9��ůt��Yfy=���V]�;����>�`�<�U��;�{3�!��w�B�<wu؛�8W��~�����?dεSa(�p2N�4�x�d��������"�� ��Q[��T�}����gH�� �pu�c�aQ\��	τg_=����5�����	̍���h@"�3�F�3�Ը�L+yDrڇ����P��n��9}���EΫ$�(u�����j�{� ��E�}��?s�C_� b��@��7���J����O��R��1#sH>3��=��0�(���>�fq,��13�T �N������� #�'�CJ��&���.���0z��F~��}7ͼ��HE�ײ�Q��i�X`ܙF=�M�vw���B:?���W�P�ذOä�lx��<{�]x%I��H?����z�q�#I��q��U�ш{i�m����#�fC�Uh�W-��~YZ1��ף� �r�I�uDm�����5ts���MfH��ä��/�D�]�N��G��,��>t>&�GiF��D�i��2���p�5��t0ێ)���τn�;�&���#a���0��=a��Y�F�6���(���	��.Ҷ\�\���1��������dc���7諢ǣ����1"��8�̇��v0������!�T
L����-�Qj��o�4�r�F>1��(>���d��`�;��A���2�h9 �8/�s���ڐ�@�-�� ݚ��nj��m���_Q�[R �F'zʹd�U��L�hl4�]��3@(�xܬ���w[~6�/�f@�62B���-:Hi=�XhY���A���WH��>'%�`�Ow���H��ڹ;���yj��ޤ�6��V4ز�Bgo�r�GՉ��
ÀѴB���M��Y(y/{V�:��B������@�J7�-��� [~��G�������Q�i�>a�(�޿��sٙ�����
���A�qb��	�$%�]9�5��R�R�T8�,��	Zđ�����˙R��x�ӯ/��|樳�.we(�,~�<\�ٛ��/~d��$�uF,�I������2��w}gA���f[���Y5��;�|��A{���@�y��"?�^����S�*�	�� �'���L~�[��H�@M�WX���~��Y<7��N]'�Ҷd�	�w���jD�ޘ�)���j_��J�i�ٚ[Gkn4�z"��[X�@~@&�j��i�^~���줕�'��\FBc	�nƈGۂ�1C��N�[1�U�����^h�yf��1��R��e��$�r�+�����LQ�&ѹ��2}�/����*�f[�i"d�M��n�ŭ�d�*t�=��	ԋ�R�/�#��� z+�ӎ�D��ֱ��7	��m�0������� $'�d�=M4�b2��EB��۫����c�	�*�)�E��JE(pA,/�	a����WBb�6Y9��m_��K����U^6GK��u�����ӌ̡�t�#o��˙���SXu�l�WTM�ȭ������ݥ�.>ٹv�n[b?��t��n�xr�K��3������ʽ��K�t��3��ќ5y�Q~��J<�R�����&�#> �^*g�)�R_|v:�W��&1&���K��D�s$9e�}��Gd6�/��R%�cË.,��:!��	����z�������Z���66�b/�8����:�/��SqŻj4��5�`��
��J�@�D��(�(��x�	���m�\�fk��_��a��	��w<����G뼈IG�B��=>?`��̕/�	~~[������Ҕ��/�I�P�q�� �"��$�a�EW$l�s~gh���K��<���e�ئ^Y����[x/���eM;����V�΀8�寧�<w�G�Y$����1{nDL��n���r���b�r��<��kJ�����������6�2�)����*�yT$J^�/��?H8���lH����"��G�����Aѕi��w�����p��ٛ����/ZX�f&J�k�s�yH ���vdc�*�%_�t&�|u���v�Е��eK�tO���J��B�M�hHL:���6�ѡW$��CIF�:q(��]ٹpF�X����G��$˨̀��Fɔ���X�^�ڷ�O���w���|�cl_��u\���M�Zi+�0��9�5�����X�����o;e����`ϐW�w�X`!��8�N�֦.����[9�Vg5�/Sr�����U>=��p�+L��~ӗD�D��������q�ڛfYm�L��3��tBg]دF�N2Ç/o��Yt�'�K��6�+�~aۍA-	��#vQ��G#d"����k~��˳�+[#T>aa�^m̈́�Xh�v���������ѻ���h�Y���oGJ�o�>�8\<�����E���z���:}���y��J��b]]�7t�~j�uGd��j�f"�>����O���S�-���c���7!6W�/�M�M��.{.�Q�b��G���g��� �#��l�0�'o�l`�|Z>�Pz���|��s��T�6����#�u�i��t��9�4��m׌��c'� "z�c=�)�[hQ��M-S���Dӝ��go���5-K �Q�"#3(j���Ȇ��`�O��~bz�z!� ���T)�f�ӄ~��[x|���3�q�x��$а^_����N���o�J0^�V[�������}����8W''M5�g0�'�����1쏞)���I��q���<�w	�0P�SzY��2ޕ�([4�׸�^��n)vᓽ�Z�7�}p�ܶ�ïh�o��Ë�A������w�StfI	�Of�2W��G�j�E[cVsPG�����[J��3�{_�����R>s��ɋ:��eD���sg�)U���s�!˰�#ky����Y��<��~wۦ����y-�s4��s赤�_[�_M�~292>�7��0&��9��f�{�"�듳��L��[�p~n�����ǽ�x�[�W��)J�F�g��m��&�@���R����)�������6��^����ɷ$0{���"��- �/bk��lN����b��X�,�q�SZ{����]�Ǯ��WF�)I�u+�-q4�5ץo٧VF��s��Q���04����D���뇱X*�#9l���i�O���ܚ-<��Z��z4�����s�?ʀFb�8���//��3�,�g���
���.>Y�`�^ a�I��:C[�{��^#�h3O��ŧ�ج��O&�[z�<깾�]#=��l����u�/��[��X���!���!�}�>�)��)�8�Tc�b�����b�(�����A.d{$��|���JaDCf��Ë��3&9k}��\��t���f�}y,42"O&0yC��B�[F���&���K��[I�gYL��_����_�֙�W�9�6�^�s#���<����R7%QD��T���t��Pd�I�����f+�)R1D$;ٷ�dϖ쳐}��3f��<�������_�y�s^�9�y�\!B�v(�Ζ�6�vWK��ԁɞ�
�1�O�wMk\ׅ��4O�Z�/,_(�в��,VR��ϧ��^���O��~����B����#�� k���ɳ��XD>�=�?�rsJ{.)=a7�R���8�X���j�l QC����R)�R ��u�iT�����DXYRT���;�_��F�ޅ�;�������7���\j����U�r|�-�f�#�_w�h	<�f%mRa�+c��SJ�/�����I��}�`��/Q �^���b����J�T�" X֕`^�ew���)[s��:ߖ���/�ǃ�<�vrO����:�� �'����3^Z�1
�E�����mmǂV_6����\��j|���yU���PoC���:�)A�� ����V��)!����$>���5�yWfϾ�c�,>�x]�t��@O���3 �� !��\��2��7S�j�d�Y>��S�D_Es���	���=%u�G��Yo�:������M♜�֖s{���%=?��R��E ĉ]���'���s7�x2`����&Dc�����a�"�$A+�m�]��<Z�}�as�6[h6)\�+�NM'�����\�@ᦕ<��^�T����Pgq��H�Y���/�3me�9��ub����;t1RY�4�{7�����bE,��n/~���!���!�9�#�4�h�����V�#��!\ߡ�ǲ\�&0of:6+�Q���J	b6����U��v�i�������+�)UN�i�\1�vR(��O�.`[E�/�$���s���jȲS{u��ԿQ�Β1���n�CA����|z�O��Ȅ�r�Nq<�L������P� �ݺ��(��u�y%, ij(��g��H�}��0N�l;��3���b�2nh:+� ���W���f~y˅�}�kr;�d�
�� C�ꌸ��f��8�L�~��ވ#��5�zՎk|�9 �Y��4��G�	�-I��BÒ�J�ф�3PU��c����'�$f_�=�.zD�B��a'W^�������v��̔�d���3r��uG&��Bֳh�D8AŒv�7��b�B�Xc��Oh(� �q�zz�_�X�� ��O*80�~4�ҮV[���D2�n�#�gD�|q�< G������.�\>03�Ȩԉp�ǲ�s@'q��Q�3h�����G�6�=�Z*��ʚ8��B��&�4T�;�[�8�м��ͧ���ȱ�c3{�UX�O�m�x�R��/@��{�[4���S������;�摪��G)�/�$�5��J�l⏠T�k�&o���c74���V��罹��U��t
���ૻ��5�IT���d+�ѫ	=�jn]�U�e.�r�2�����%����i�O�����ms� l����?�7ڲ�X�'K�>��W�{)�Dv��)u3P���^�A��Dh �c�����?Z��;����}���r�@y��X�&?ي�
WE��7hrİx����%��S���n����i],0�4X�t��re�i嚫��ָD��ʕX{��95�*�H�Ɛ�h�dO{���^��5�ĳ�����;9Q?�W>��*Ί�l��2��IE�8y:�M��Q�jU��������I�y�<���zX\�b;)�]^�;��b:�|V�%h���@�g={z�}�/�C�c,�����g��Qaw�" e��5{��͛�I��S���B����HɛN%UK4�@�����AO/ru9f"2�ψ2�}g�
��h�n�<l��N<�>�K�I_2X2�J�F�T���@�W�:U�$9ܪ�M��4���y�����U2��	��H�}d[�A�蟾�͹2b�%�.�������!���!�=�P���P��2}>(�ZM�\4@�����}��k�Ϩ���&t�o[����SL�h�%��Q��W)	41���ݳD��%	[〉1�I&:+�O�	�{(��X�33<��`�I8�Yx���R���0
!��pQURĐ��f6%s�h��@R<��b�P���_����;<�1��|��o��^��z�w�F+B����~^�f�'�Qi�����(���o��Wt�"��N�
p�e�\��������u]�v����ɋ;�r��t�{�#��r
b���a<�.ݩƹ&��<LDl���3#�Q�����e�I@veʒb*ǁƏOF��Z�t=�ƥL�_GEs4�k��]H��Ǵ���9ݯ�1	)���}P��9�V�|�`�Pm��vS�#����@�N�!�yH��Oם��7��/� +���㶬|�}p��
�5�WF���mg�J��R6hIH�����8֓����yqu]`D쇚xgD�z�64.AE��,8����3P2�;IX�����;[��:�	̦�@��v?&�~>�vKxD�8����=aA��Cm�� �'����]-ڸE�q���"sA�Z���g��V�cv���O���s{��I?H���'��82�2��~o牍Ev��VwmҥA"�)ԣVJk���Q���g��c�ܐ�B������I��=S�C���@��c������q|��J���z��n��zG�'ڻi=�q{� !^�B�j����՝x�u��ߴϔLp?Q���r���d��;7��n����s����:	�1�	(2�'�E�O�?����7�:��uQG�y&Y@���]��F��+�ю��t'~��f6��SR �[� x���;��x�$[ڝ.��͙��!Y�(ǔؼ��;�,)@V`7�O|�]m�ub�'f�)������'ߙ����� ]�����U�X�����
k�M5�wz�xh8��v(�r�=�p3��W����`]�@��:���KxW�zu����q�@�2����Fj��}���GP�
i#ϴF}l�t�:d�{��� ��PR��/@��ˑC�I˄$w>��"�
��&���xu�������<T���6�~�l\j�����v���������7<�.5f�)��c���/�͸O5��	\y�V����4��5_E@h�W�G��=�ȯ��gc�AP׈��"?��Z2}ZΏ#��4e�td�С@�f3@˒���*в٤?L���?U���s[%���l��\)�˨M��g�&7��*)���t���o:J|����A�D���qj���`L���4&���J+/�9A���`�%�e'`e9*�i���։��NH�\�\�W"�iӬ+΁[@��[�iY}}
;����� ~>����W]z�4�p�2�؄��C�:�����=�W��Zn���,J�]��W�������Tt�v6�#$�.a���/��r:���jպ?"l>{/EL
�AK��\АR���%@��k� PC ?��`e�n�PE�.B;���>*i�G��7����P�@�6�j�A}��;\�xq�r�_*MW]v�j�ȟ�g	fF��?��|L����ߠ �.���5���V4�^��u$N�MM(I@>q(�x�d�P<Ю�ϛ�so�U�ۖM���l�qM_e	�g�XL��q�*H,���=��ϣ.���B���:T-���<�pj�*D x^�79�χ�ε��W7�k_Z��n�1$�pRjS$�� ��oau�w��P�|����n���*��ó�8����B�4��i1�{���o�B��}~�Wܥ���������**�6�	�o�a�9,�zZu8�:F�u:���>h����]�\��O�Yih�4RZ���S���S��,ޘ�/���>,|�6@��ɋ�c�p����=�x=�;@�����3�|�=3��랠V��{���������0
n�x�
��
�e�"[_�������%���ߢ*-l,��@u�������(�=�2�a����[��6vhxh�P��p�q��CRC�2��#7DN���E�QV��o�����x����l�C�W���"d���@�9�ㆁA3�2��4���y^��@tG��H��'���C��@#}6�T2jt�mh�МS�O!C��޷�,��ing[`k��Gj~/�	�[�$Xs�|��x)��c=�GB$*�hX��ѱ������lE�����q�@�b�wVs�^O����"P�}A�)��3��;Ra9���w��1ͷ�T=��A����n�j����\e���Es�
�ҽ>��6���?�0�p�?�6�>�j¸�r�H���S��j��rF���@`�77���V�l�-�+h�إWdj���6� ���a�%� �%�i1�$��nJ�',OO ۺv�� 6� ��#�_�{F���ފ��y`��fOA�ٔ���Cf����fx�,�Xu��)���v� ֍��z�x��̙�[��[��VwS�_"�i/$5PG����7�Ҋ�P����f@ӀŦ�C�P�����T�҇����Y��)%��-�˵���v��R.�O�a�ˆg�tj��DJ}H0Nk</NI9�a���'�h�6@�a��xQ���)�$^���
��:�?��[�!0�����\Qg4�CX�
���x���
��y
����p�o�$ӻ��0�ة��p{/3A��������.����--��w��u'Bu*��5Җ�m�� }��kio�]��ʺ~��0U/r��(2\pPzA|������){������<��d/!S�tС�Cm���$
���ܣ���!v��f�#Ûo����M�����e�4�\{ �A�)�����}�P���T! �9��J���OEG�ʭv�;ϳ��k'5�9�1�+�D�a��C���&�	4j$|b\IK�8���y�Ԅ���)t׭��!R�7t�c��O51o�l ����3߻�P����G�42|�ye3��@�1ʽb���(vK5	m~[Oc�"٨���[#��D*J �"�h$��Q��l� �U
��Khxp�'��4��T�{�v�o�X@��Z1�F5��l{���	�g�3a���k��C>��5�Ng���&��i����ģ����+�@�GH�Ym��jt�$��*u'��t�> ��h��m^|JשCٽ n�*#G�\_X���ɝ�(�8O�Q���`�Q�X�a���|�-q:�ku(��������~���/,��=j����Q��Ts�L�aef��d�;Xל�g��yE��+�SE�sV���do`=#u[l{��r�~6?�u��`�8L�>}M;��7��_�Q��y51�?qX���*��A�B����!�S܁�v!�jx�h�m�2�;�l��x ^ �6| 9����x6�p�����@�R�٢�w�:Ō{�pK���4�ԂO����R��ii?o�;�L��CxO���o(��S��H��&AǱg�3�w��eMI�O	�k��$���O�I#���f�	�s3�NU���3a�"
�sr�qU�oKܴZ4s����_��6��n�c!����������4�V�}�k�F	6Rq��Q�8���J����~��O6��� �~EF螸��>�D��+�吐AeTq0��FX��
5g>֞b��i�f�ii�5�II�E����.����9]��&�0�;���(�G�oB.���C��\�+z��w�tL�G雧%?w��}�7�E�n��Z�fc�������CQ<b�Źs��5�;Q���)���-��J68�O�]�f�E.�U�ᛣa�a�}����R��\��I��YS�U��߆��ޔ�U �䴒2�\���VٟQ���
����Bl&��Il�w�݅
���JI����}O�O�jQ��G�%������=g��~�JpRA�L�i3�N�M,U�Q��/�\�ov�t�hfS�C,�����[%�TnUE���p�u�m�O.��s�]Y^�ڼZg�)����V�>I�]�7G4�F��P�����A��oÆ�p�����C;�.���T��x�|I��ν6p4pA` �>8`�m����!�.�,ՊE��9<�� �Q�M ��\�I�W�q�$}��;n/��	�"�|�e��2c/�CYo�����uN�,TO[�^\�S�\�}E
�u\%���^�.ª�M껨�Φ_.�*jF�P��/� ���C����$W�N����YH���>�\Kc��a�V;5���\�5��0�����X����������chj��E�6�N܋ E���Wp<��%�K8�3]��OKr�M�g��T�����"FK�w���Iqmsu���n�8�\Qš�-<b7ƃ`�K`�̙����Z�Z=�����U��u�F� Θ�#b}�KLY��±�/J�nH�և��}��[&�w�+G:q�%-j��B�	.�1_����6U��s�}X��ϟ��ș�Z�������sm��#�J��iH�֖2�4�<ɫ��ˋT��ZG�PӆO�����A�t�:����� R��s�}�(�z��<ϗ� �y���%��@�7=��6$&�B�^C�2���������mJ��yLb�DQ��|���5r�?5��VT��}ec�)��,
�S��Q3?W?���͘��Ӕ�Ǌ�Fj�𲡋��l�����)r���b������5M��o����z��7H��ٝ:�AB�C���a���g��O��N��~����pY--��~K��G V�<4�j���7g�F�eZ�,z�� .��:\\�g����P���X�Gi�1^ЍƗW�L�������:P��]��!���2�����ȡ�<��=o�������5G��ҁ� �
y{�~��ҿ@讥����#,q��Q���4_T�!j�G:f[�/{�)��v�}Dc��1
G�����w�_�;����j
VB�5��HT�Q��1����^,-t4}���=�^�i'Xly[���ף�S�:��^P��������i��Tv g#ⅢNq��N�x�{n�!�d�;��?�c_��3��(�Vޅ�}ӊ�]I� }��M����`�+��2F1U�#Ԓ��5]M���~iE�K�p�J��<y1&<<q���!����O*\~n<3��~n-�m�3�,k�@�e���8��%�B�n���8��p���an�V��d�pš��c����q6q�4��	}��,殺�-�)�/�� ������߅�מ�M]��n7���W �i�4�:��RB�q�lK�·�Sb�}*�n]�Ib��0T輁a=[L9����h��fF�o��5���۾$L�=���S��<g��ؿ|W
1��΀3�%0�F�������G��V6:R]�w��\r��޿$����_���
3�A?&��EQ5�����>օt��ofF(�;؊�JԞ׊�sS[y�/���ˡ[�x`�~j�7T8xB�\���C��잜�0w�t�`��p7�]��*��O���&��O�u0�\7������PY��B�r>푁Q{}c7wA�.�4��!�������y����j+�h�۟x�s��|t�;+9pxc�,��T���� ���\�m�	��G8~'@2f���F�A^���4}�{���m�X�L\)��l�S�k־|
b~{;���/�c]8i�4���-�/�<�9��W���~A\X��ߎ�}��������6}�uzz��I>
em�L|�w'7P��;U�EV�-|�m��?`��A%��v����I�?H\`h��o�{�ݔ�V������{��|9�2���_�l�ՌT/g�-��6�o0@njC������F�`��No�kSU �������P�,���l�%jG,��[+����RkĒ,ga���!�������1���z�Kd�� �i��#�vS��P(������}N����Z |!�E��\���SI�k��|���?�)>H�4�"q�>/\����(��9(rthw�p��%Ay��y�W���ny?��&p(������+�׍�1�Ν�!Uf���g<R�h��	v����<"&M���?31�{��~I;�}�ѡ⧨��Kr�6I�0��q/����2�d�[]1YY��3�؁]ZDP�d~�6Ū�hN)K'�a[����
����V	��3n�JouTo�$::����N����5L'r��-�`�ڝsm:@ld��h�{I�"vJ?Z���m�DT�.,?
���_���/`�씦���o���, f�gg�y7���SF�j���*�l�r�66Phyf��5���<���@ø%�h�u~p���z�f�4P��?�c7X�e�|��CVw��G��O���+�y�?WȾޔ�]]��f��� ���F
0�1���z�:-j�����S�~�U�҆��/劃{� ֖X[�Lc�<�jb�s��FH��̿�/5�?��( Z��p��4���-���L�o��� ��"�?-Q�(y�����{�NXcunc��8������b�t��D
BHY'�PJ����߫9!k �m�Ԝs�%�q_�Wm*\�o�i'���7���
1��Loi��-M�����Z�t�Ȯ�2%t�J_ �%kذ���΋���G�.7��S�FV�\�`��׺�R��qM	�zI�қ���~�Mu\��~K&)Z�m�,-ψB�Ґ��R��_s�%���v���_�c�wX���q�i|J�r3�~f����D�r����l3	<�}�]u]MZV��h�����?�>#2��n)���$����5���į�{ye8�:/̳�3���t��ܻ�(�.T4�>2,�$�6�ͬ�w�#ߔ4��Υ���z���d������>�]��_s�3��� ��(Y}kJb�]�ߪ��N���L8���U�d�K��q^+�C7v�=\����^+l�X(n:�Ͷfw���+C3��\���]���߸,`������,Ҋ�!��WQ��B���G��c��=���Ш���ŷO.'/c�J7��Ԭ�������j��ԭ��R5m7A�>�@��M9����цjk]���N���W*aP��% S� �Nx ;�G�gw>�>����y�p{[�!���!��ပ�WOz,�(�T;
���vv���dI�V&"q9�86Um�թ�9�ϣ�O��y��j�R�w�A����_�w`�a��:���g�� �s�nx6����9���jF��l`�_)��
���\>�ߠݯzu���+
���=��j=��8jg@�Z�ۀ1��;����f=xD�CV�G��R}�1��oK����A^�ܷݔ������5f�f�~n(�`�kT�3ս�4l���vR�sX��/�i����<����Ԁ{����	6/�o�����2���,�țwhM�?��<�,�}��=�*�B�Nds����È��5� ?�N�l��ǑO���)l@1���/@�>/�E5��+�Q�ʬP]XO^��?�#�V�d���Ke��:�,@`�0b~Iخ7�[UrA{d~/Z�㋟��s�	�%��
�0� ���S���x;�����_��$���{&���r�|������z@�����^ؔ�{T�Ko���ʦ7�`�{{�}ox��ϡ��=�0�|���2�z��9�;q�_C��.��HZ�RU�X�v�IgU�؉_��	��i��������+=�?���Ud/΁G<�F�6��FJ�-��WR����?\�<�:A׷���6{�I��h��nOߺ�y�9�N�k��uv0����-C��^�2NXy���P�ls~�r���Oxx3���^p�����cl�d��<ĬeH|�V��0���=��	yX���!v�p*[]<��u(�=�����u�'p��%�o�Xko�q~N4����oI�)�u��>o�����w��7/$毓j����!5-�+hP9�8���<�� 	�<����@�Ojy!��գ�Z�Fվ�ZZ{��0��]��YH�L4�K�+����)k�o9��Ԛ�h�;b	Ɏ9X��;8/4~5�����i����&�`9C��������YW>ffda�M���V�7I�`1�H	�x��	c��� �!����	��?g�֮.��h����h�,��z��{&�͌/8	�y:]�3W�`��GwR��)gؼ��:�b���GdG6�$��1u��jR�7�-�X� �rk�iŀo�kt Ӳ@��OS�-~Ҥ����rZ�2�]w�f^@�E�!�^q@@>��}.�It����ԝPT������@�M��/K�V�2J��s݇=�cN|�́t�7]�U��n���:��إ�}�rn����0�qm����=@�i���z�QV�� ,�i���R��r�d"�8J�*�x�.sDR�hŤ�a��;8x\�'���8��>wWm�Dy�R�&��|c?!�,�Mn������E�ض�`����b�-L�
uq�z����g��)a3���UZ�=(x�g-���u�x�)n��D�I2���}�4�[������y�?�ȋC�>\
C��g8����,W
>�t� ݩϬ���~2@�<�&vX�Tf�^��N�`�@�d�
$[�����s�X� ��;v�=�s^�#�+$��G��\�U@M[�B��1��� ƅL���&�%ʐ�g���d��c�o��P�2;k��'8�G�+���]��T��)��n9��ڐ����[3Q��,����0l*\Adb����h���5��[N��|��SC!�8���V�/��Xx�����'ކ��/�U�2'���2����~��AeL�R���/��}վ2�����@!��z�૩���9P.��j�#���*��������j��lۍ'�Ȟ^���ʃ������d5ۅ�/��̦mg�+:��~�y�S|��=*.�FM묖����,��!��������M�Z�唭�ޱ��g�J�~eۅ��̥x`R�J̡����:%��s��1w��؅p�e�}[����p��{���@MM���D_cM����#�$�M%��ʲo�m�L�uA0p��m������c|7��<�\���r򞩮]�b��$6��ۢ
�����ZuSqzr�Y��	�A��W{K ����լ���sx�1 z�ǫ�������I!��7�/0�*�ت��mguϻ8[}K�L����O
�<ɟ��I�n�aU.�s�$����m�z���ک�����:�q_J��̗��8�����<�?l��g�a6��Wj	��7�'���z�謵�V܅��>�;��n�Ĕ�����{e�$��c�K'((�ɢ������m�*�և�c�2G8�}:���H2-�H���.nj����ܙ��Ofo�]Z�b {�[Jr͓sjK��"��׮�O|#bE����e���]���]�=���B�	�0��$�J����Y�����̙�j�c�X�aN��yX�=�A�p0��z:O&�mr�z�]��kewi����-z�Y�=绹1g\l�v1��*U�J*��d~r��\�����]��|J�Ne%�k3-�T����t?�և��-�˙�1m�u(4.�C���f!IQ�4�N���~;H���no�0�/f�l�t�n*d!W���OR��eYq15�~~]��V{��y�,�Wȷ����6��w���=|h���V��B��Q�D��[�c���$m�*(���i���5tG��ť'퇻���b�\�:ۥ��$�$���>���]l�R� C���P�#;zf�`j�@�K�J����$v(P�Ӥ�ec��M�X�,�}X�)@���V��*�����}���<���I�K�QUxj���=b1 �R܇>RO�������	~$�"�=o�CT���F����� �����}�������n� �U�� ����4P��<�H�C��|J�E��z��;��dq�Q'�P>�a�q����&b���ߺ��m�>� �T��r�YZ7�_��c���ɀesaiKX*�Z�2�W��\<X�K�|�[5��hA�kHp�4Λ[�ٙ\����K�~4>w�Uv�^��0�Գ'�X��c�p��GA��H5���G��ځ&�h�s^�\�G�1m!� Q��j�u�%u�f���yi��H�EV�~h�q�8X����X�؈�fpH��u-�|5��+���nP(T�T[y�cxqG����ωS�^-W4FJpc7�9�1�����xu��Ǌҙ6��G�p�T�a���9X�W{���$����vo�zs�zx����)P a�έAC���+�@b��F�i����y��w 2��K��z�D� =WE@l���#���4pe���
�P$% �F ����;��p�e��ʓ6��;V"{;1W0����$&Fzk��Ĭ���o<���e�`�򱂑�:��&�p}[/��Sbsn�4�u̐���EFH5Q"T�N؅���3�?�Qcl���A'Xt��H��$kV��"U�G����W���ݼ{v`�R8(lŭ3��%c$��eH�P��x�`{��λ|�H3MJ�=�~�.\t����R�e4�4��e
1T=�����i�B�[�E���e:�1��H�ȟ����Lq�upR�-!�<x޻��x�����U�w�<`Y�����!5�vCx+.�I�_�����̈� � ~ǭ��ndg��^EV8�͘V�T�~���)<Pq��p1���c�|qO��A�?�A����[�ŭ��T��Y���I���K5ȴ7�_��C'6��^ޘj	�Ul��[S�T0&h�=�U���0?��,[�6�/��H����1��/N%��s+�~Ni�W������X��7�U���Ej~oZ�P��Ф��,��b#�(�q� �s���ã+32��>��قe�Q�į{����w�ݑ�o��#'Z.��~��Jh�R��̓:yӫ_�4u�ټHÕ�e�MU�'ͼMR�Ԓ�0�rGT֧ߺ���1�K�-�R�ܼP����.�F�ĭEZԱ�[�ל����q�W���}�OY�Y�H�6�I.�>���#}_+!��^�W��E�qq����L>V��_<"��J���?w������+�x��i}�sP�i<�'ȟ����������.9���iC�>"��[�ދZ��X\�+���?���0:�#@I��;�f�X�Ԯ�a�r&Nkɷ��F�D{Ֆ�na�ar�WP�X,�JT�顰�Y�) ;�8�crz�H�J������y������XHQ������20�1&�3��v��H�Ģ���O��@ 䧀Tqة}+�բ�3ϖ�ze� Ӗ*i�/��e���c/I�)Vg�&��L���Rvj"�� 0�Ƚ =Ǚh�����V��jP�QWY�	3��Ϛ]Z�g�����;ws^B�)J�gʕ�v�К�{���u�',h=Gm�״bG�RY2�+�]p�3eGg�J����}|��7m���gGͧ���ڝK�ؙ�o�%�
���fI 3��9�P�p�� 5�9a�T�����%�߭�~����y��Ì
j�e����zo������xN��tU�!���	z�B"���z�䴖��DX��>=�I�����s��02����ٿƁ:�����#da�ջ��S׻	o�,_!���j}z4)i 4�<��>Rei��2	F9���L����)m3&�=��vsP=9�]���d�\�6pO�L�g*aݿ�J�&�J?����D�x��Z��d��Y�b#q��
�L�������54��uv�^jSjb5�)!�*8u����de�M��L�痊NQ��8�T��J0*>t�����;y����Y�RF��&&���������{S3C�7	��N�}Փ Cl����!�w������D��⭣s����w?�vŨ�p����_����=ѯqEANh��p�˘I�`Ԃt����Q�{�};���A/��5�eTBc�Ă�qk;T#'T+��ƶ����m��9١Jz��r�$�#��ܵ�ǎ��׸�?E���q^�j���,q���Y�?��c������@�P��i�vTݯ����]"�����R{���Hɒ0�y|2s���y3�TЩ����9�g�2�s�.1�?U!���o� �)S��9�GD��`Ǧ��Rgu�wl��ρ��-(�mw�����)��DP~J����h�c�3�U�L�{Փ�nhTK�q�K,��2˫Q��������c� p�[BŌ�o�D����%3Gʼ��Y˷�Fo�K� H�ޭ{�#4���D�vz���ըa���|ٜ��(�����JbC`ay��rL��(GB�>H�c�� �SV��U�R�
���ß'�Y<{����΀O���6&׻��Ӆ�Qbnb��w���,Nƅ98G����5��T� _?Y�9�qM��oٰ��R0W��VW7� H���RA�����o�S�~�Ο����g��x�^KY�����N��0�~h/����0¼�ْw���=����|uD�>�Ⴖ2T�&pQ�HJ�dt�T���)<e��b1V��u_8� A%�R�V�?��,~�v�#�pe<���Oʺ���/{�}}1�9���u��ֶbBf���3Y���bK#g�"�s�k4��o^�A� ���&�>:�=�	��U&X�����5c*�Veb�`	�Hڼ�K�n��@��|D��+�똑���������Zyy�t,�*U��p%���p?X�"?�(�?`M�A�~h�#���E�?X��LJ�MI��Jг|���JeA���Fb��|����6*�DNefż ^Y[ՁGc
��`��KV���,91�E0@0�]Æ�R�MU�H�|@��Eo��$��~g��}sp3�XY���kE��t�%o��	x4=�Z\�h����@���S�XK��^5���2j*Ɍ����С��_����B��!��J��D�n���@u!���Nּ9z|>���&M�u����0-}�����z���p�&��Z�P����*Լog��s��e6�\�����H]�CX�~�.��L����ȼ�g�n2�ﻖ�Qnh�Ժt&�.�qh5@ �_���Q4�����3Q�O��1�
����p#f㏹��\4��Tc%�0F�>�%�\�)YI��q�^[L��5�EG��֎���C�w�(��;Kl�����ɖ鷛�qo"����v
J�C���F.y?QB�X�^؎��:ή[`h����<4x�P�Φ�<&&�yI�[S��/aJo��OiE�QTb�L\V��{rG��|�����9�� �	4����vCW�J��,1�}�JUp{q�7�M�%�u��Ҏj��L���=�B��(���z9�y��{C�9�j)D�=��/m�F�G���/�;�x<����&���Į�I���lbQ�0�r�*Wŝ��<�\0��VX��Q��g9Ce�-
ì
m����T˄���FC����EZY@�����;+/�y(��N��&�&3d�8?�2�ȅ*�_��%�'N�	B4�|)� Ii��
;j��,��̨��}:�08��ܙޟ�7�G)��`jMll��'�[;��C�S&3U�;��n\��2�G�8+<����b>���4�j{�	�"�݊��37oٖ'j�C���^o�)���nb�Q���2(�����U6�W��e��i��89qF��I�5�E���.��P/=�P��Ul�x�J��t���hD�X�EN���>�ș���\�WXۇk�~:�{Zc����tC9c������K��5���N�C� �(:P8A���(�R~��	6��Oy!-�3�(����9#dB�F�D�v�s�`��A�Ml��VX�'~��F
N�D��M�����J�v��ES���/��z���EmpnмP��O�Xm/X��jd���MFKgv+Οiڛ�^K�N{\EӉ�*;5N��Ti_�d�
�E���ݜ�Z��>�\��=uP�Կ���f5�,<�K��q(���9�W��8'�*���{N;�>�wb��>�m�ρW�X�4�j��/��i�ݽ�$�V�k�j}�oʞ��n��WM�+��m�.M����V����@��4a�@�fv��6	���0��*��/�|��z��3���YCP�@h���]�cyd?�����;E��rA��3�E��1p���s�����G����� �'�L� ���j ����0�}�x�O��`I�����a�ʿw��B@�U�`�;��ԃL̘�z�����OT�d��%>2Y�m�>ۏ��h*"f\�����x�����5�GH�aS<��{˽��Qd�H[Ţj��OW	vU��������5z�o=&���:`�*�}5z���Z
삥r0W�0�l�D�I�*}�ueT��4��[mI;�	����Uʲ� �FT�(�a�G�iS+��_���! �Z��� )J�)�%?*
ީa��cX�D0��G��r��f��r�*x�&}�>��`ٺ(m��R����}8�`�O�`\��dSLn������pY�]9Q,P9�g�
��~Sy�ls�y����p؋�Ŏn� ���FhC�F$��433��cx|4���YY"��jq�L� 0��a?� _�V�>p���v��݋lv���d2/�����юq���Kb�a��>KܸƆ@-����~RZ����?��&x:I��F��5�^��ES<�|����Үt�:%������
�@�dEY��G���ܜ�]�U�k�p2�k���02��Srk�릢��!|��mYz ���M���Z>Y�jMd���2���L@-O5l|,?�P�G09HB���^�fب���ax�(ٌ�����Ոb��2I�G��ӨƉ��Y�ԁP~���e_Oz2��Ѐ����^�h���ˊ����Q�7jj�h'8C�7�h�������̼l�����٨�7��_�r]O|ǉw�w�*o�s����ߣ���3�4G�Ź��p[��?��g=��%i��Ě0��y����F��
&h=��`����g9��[P�����2N�Rn�	*�ʙ��f��	,F)�a>�XUg4[��PJշ���FY�qvX >#&VS����k��T�<�N�!��ɂ�y.�ubO6�P%:�A)&6���]y��. �}��q<��R�o-E���F���ҟ�>�F���<8|�7 7:9���o�ǰz�,W�ѹ�>k&mQe\J�ѝ��D�ЈcC���6TeL�'g�}[�(\	s�c��"Ȝ�����Uڒ�`��c�y��ʂ{r[t˥̾��&c` �VIL�x���Fh�������2�:m���q�N��R�Ȍ�^B5�1��E�G�~��&}�3��}����Wțe>�V�]��A�/���ˊT}R�J2Z�o��c����[SÏ�b=���=�
�~��}�,�z��f����i�CbnSw���S�������)�e���a��NZ�K�ϤI�E�ĉ�O�)�؊�2��� �xo&��Hހ�:�2���z�غD�lN�m���:,���l�2#R�C�eS�`�����WLJ�d]᫵[U��4i�����QQeY�p9N��"H�-((ݠ`�
J��A��`���%��((��
P�@@�H����
I%�P�(�=�ܺ83��������Y�캧�N�~�ާnյI8��!�A��J����"��~R1I�솜�w�|�b!�����L�D�t���z�L.=YW�3�|����q�O�B͚o{��J����y7ﲛeV��V�1��p�g���]�\[�u��l��jƝ��ؐ�"��>;��R��sb%P{;���6:@�D�>�*|v���Ws����|9�S�fBMz�
g͎������Ǐw����M�FȯKm}���ۙ����b<���[K�e~�l�@��MZ�[�R�B�`]�j�Ǩ�&���aA��5U����"�@o\r���'���|ˋ,_�9�/F@C'�:S��uG�������1�LT���/��б*���NN+�Ӛ��W/"b"L� �aP��Z*��ƀϘ�D��K��1>����m���_�o\��`�ᣩ��"Y��x5� ؄���j7��|��~R���rF�l���`�rwJٛu�)%�W�|fS��e긠M?R���+)\lST��v����xh��.�K��:�s�B'�x�����LVS�cL��|�#	�e�
��WfWz��ښ��di�}�Xaz��˸�AT�X����<\����xY@Y����.����+���f4��Dwd9{�����a����m���<��B�󄴧�gظ��+�/o���MԢs1����R�
�t��v�x��naU(�'#"9�3�=~u"����}#��CQ�C򩣔��"фn��ya_�Q�2�Ⴡ���"�!��:��z����+g롻��vY�J>���9[#$���}rB��}�E�n�F7&�;��+�<u�p�3t��z����%#���j�g�q�R�p�ͳ!�����k�/s��w5���n�io�'z���6���������5fg�К��慬�Z�{҅�4w���/��)�>n�D&�����kG^֏��,����poI�����M�v�?XM�r?��:����4j���jw3�m�m�qeN��zy�4F���U�"0?(���	�s�v<��,l�q 1�)HQ'ݬt}V�t�8�`Ej�_���	�yq�
Œ��= T������4<ߔ�E>+�e��5h:��j���."ty�k���{�qrs���'ݭ<]������0�),����gh�Qn��"
���zw�m��R[���F���*v��8��k������Gr^�D�ls
Wy��y��^Qp�cX�5h�c}�����p���u�����Y��;��9P(�/�)w*�G��1�'���f�H����8�kj��(���i��*�ӏ[z�DLz#4e#��S���@��Ͼ����:]c�Zg�h�0׾D�"�h��z��W��w���R4UN�)�1��i#���Ҁ������CEe��NJ;�0��A�6��E��zW>�\��Z�#mU�&�k��̳�v�fҳ��0^�p�q��lKp��9:���,ȭ8OH#Fπ��U�<㧥��a��S�^yu�F9�2���u�;��F�һۣ� �$6���������͍mor|�{�P�c��3��S��x�b.uc��~-�iq�]�Bd���]�����ՀJT�꼀���pM��pi�'�+/fl��}��l���� ���Qv��-�j�Y�(F�6x�Dz���!�	\��n[�ݓ�%�q=�B��Ḟa��_ ��nμ+^.7[����W�u?��c
�b���c%astPv�7�e��5UgT���'�����,�G���^�ͯϳ?}/�W�B	u�ݸ��M�~2�"�3���]�����	�>�+���sz~�*��2���+����1}:�N�䩛��YgX�̌�`�u�˼@&�{g?�0�����:7��A�Z���bwa2�E�B�ʂj������\��
�a�B�cF������=��=ν��Eh-�ܞ]��M8��t>h��ʼ�њ<��;>�|�X�T�f���h������`��~��צ�L��.�9my��5�'�֠����E�<k\(q�h������w��Jc��_`n��Z�)5['�>���¼�lwƳ�Z��2u����Y�~��1��=�S�ݒQ6�Q�{�0׵=�\'� �[�r<��-�F�5�o��f˟_|%P*���#O�P#����HѴ�ò�����wҰst�W�w�0�E�(�y�W��%�U?����J�Z�]��˅�.wݰ݋������)*�Z,M.|�����m�]��ȓV���*�!%�n
�
���s�P�HF�9>lwxc!�:,�v�}8{{q�FżZ��F��,� ?�L0�ȵ�҇���G�%N��8C���M]�Y�����\qo���8�r�u:���4����X���.�"�6 ���'΢-�����`�T�A M�~�z�U4o)U9���CP�$��3*Sx��YO6Ep����.���7�j�y:��U�+ZT��gTs��|	R�NNЉ�Ivr�є�ީ�4F���eV
�����C�
�%���u��z=^H����C�����Nkj�
����f��aa�g��`�܉�k��:Hq��5�mϰ���	��ڱ�	����!�X� ��:�x��@���ʹn�u4]l	r�xz���o�g��%cx;���.�(�NG�F@��������4�I��tIy�hW��`[>#l��@P#t��&;Y�
j�k�9ۍ��������Zt��`���k����:�D���m:Ʉ�*��̲7�d�6On�P����#T8`�L�j�P�V(�]�#��;�g��aq�SQ���7q;�I�����q\ͭ�Z�~`X>$���6!�m=5�_�2%u����znW����@��e����Z�_K����%�sD��Mn`5NF���I�*v�O���t����)O�z�η�/c�������8����5�������X��-�쇍i���u��M�8%��Ɋ������s<�Π��p�} �,� ��mU�Zâ�  5���6�V�5��("0nElJ���(b꾾�_[��Z���;�ɢR?�C`͡p�SC�92�&:N�D�Z)�,2�AL�b�k��Y0��4a����g�ݐ�5��o-$)�^�GjB�e��Nmw���%�-��IX�.�DL(e�~�����s
>d��&�m9�RpFG�ܼ���|'�iv�Q�B_��C��L�N�_OS�-p�zd������P��`{`�s1�4�9�Qǎ��Ԑ�t�#��c�GF�g'���gG�u��}�<���]^b�=�3��{�����[XwGYz��b/=���I/�t�䡝�"��L}���%i�ߔ}�����Pxw�}��^X����'��E-&C
Ղ5�܅�����dY���.������ݗ��^�oـi!�����Ӗ��\r�;��!.�0����f��|"h�k�����h����\��,s���:��n/vʱ<�k��X\c^6s�m�9��������sH¾��7<,~/�M�� B�ܘ;3�$~�z�M��?l�����;z@ӑ3J�l];Th�>xC#a��g�9�[`k�kZ�<ǹ�N+��}j����k��[���=�,�ry\}p���H���(c���Jx��y<d�wa��I��ɸC��]��Z��o+�ο4�y��d�<�Z{���t<�Nmi'�c	��GU]2�I��Ȥ�����}:�����sA�Ōk��W��Ż�"_|n�����X�6Ӻ�e)�*�
����^2a[�8�P�$E�kh͞}r��Ǚ|qqw��8�ӑ��oP�qz�u�&m�]��-�Ƙ����"��7���R�I�5���y�ft��ΡО���,v?�9Ğ����.�q:��1x�Ξ�/+�1�$@���}����ڧ�B8Xٱ��1�����A���z�`�t��}`�&����84zMa���p�h!�����@9^q��Y2���V���}�@��'4f��>o���@����^��#x2_�AN���RT�e�^4��7a�]i��i�C�{Dx2�|������U��z���	�N��,�N�4��	�:��9Y�umo�ƪ>�w?��	�v�}{j��1Z�!��ׯI�~��P�C��^
z9�|���������)�e.!J�i�)�G�ŉ�X �7* ��a֪ajA������U�<�џZ�߃�a���J�w���/�Ã���5��NKr�Y��>��]���AKz��W'+�Ѻ+;�����c�b��@�~��k�1q�(�|P���1b��'Z�k�:V�;�6������.7� �T.�\4Q"����	�)��J�� ���j��\����]Rh���KĜV���Q=۞�uKiK����D����`��B�=�$Y6�:�)���c>�s$*, ���@����C�[�kc9���3�zP?� ����>IX�Wj?{?3|�n���ʶ���I�D�����e�ƿ�����5
�u�t�;��Y8B�q��Z@;��_n�M�l�B;iHϛ6�g۫� �������S??�����Hf~������\G=���ю�b�)�耲�E_���?��d}i.o0~��C<�̀���s9�/�-����-��K�u��*(>ة�?���k�nv�@�ځ0��u7��p�F[n`������k�_ƃ^k{4.?o-������@����6�1um*�˫�_�M̹Г	S�؎<z��3���r�Z�5�·DLt�DT�꥟c^�i�=m)�"����>0���J,̕�a�+;�ڇ�k%5��M��( S2�����]b��.8����iv�+?�~��NKI���[��}�|-��P~���=������S=y�o�����<F;i!�����n���$dk�u�3w$x�/��Gئ�8��U%����؝f��������h A#2a�O�O�,����=my�����B���M�g�-�?��#-��F�fꎃ�9��3�𖻔=���1+��A8ᑠU7�(���=f��Vg��K2Js�;
>����:��EO����`�fm�vD�t���u��a����x+�iԎ�9)����՛ﻔ�n��0i\7=�$r� ��x8]��v�l�ů���DHw�c�Q*�VW�Xd�1h��s.�(8~�0�ԯM(�tK�Hn&�\Je�_̸�8v3/X��i�_V'ҫ���&	Y����6��ՎNWqe�:-[Kr��lC���#���U�;�:��\g6r���]�,��IX4Z�w�����3�g������Ŀ��{^�.����"�*����!�V�����ڜ��9�%����+�C��xv&�H������yq��\�e��n_�=���]+��6ފn��$k�̭��5L��={�����
�����on�O,�ۗ��O�,֍����w+����sRC��,T1����Gqe�P��ç��x��7�e�W�s�x𾯚$L�D���W������e":P��0_}t���Kk�c�VT�~%����[|+��*-0@O�2z�D�p����>�\���o^�Y�d��_�xsq����^��?[�Yӳ[���)R�������^����+�EG5�UJ�@O��@\]]�^�f�$'g�"��(���D��F���
��7'2c���O�N��{���+���y�����|&	o:��Gχ"6%h���7��]�ǁI���t�ʸ�s0���;�|]�eT]h�h���;0���|i���쎱��r��ݾ6[�������מ���ү��k��7?ؙ�^�zc��Μ���"��:�9V����M������کo�rq��f7븓��եz���~�����dwXk���èSB�)l�h9��a�3Jc�r
7���;�o��w�8������%�z���+{�'���C꩏/���$ǫ�����\+�} �x}:�n��i�?R����������È�=ն�J���ӣ~��Y�+�_��Ƹ�U_;`���.�Jѽ&���n5��U�Gf�,^��L0�5�
��)p]��1A%�+!���k�Y�����7�-�;-���Łm&����LwJC��[#[v����h�R@��߉���R�_��k��u(1�����m�Qe�A`�Wz��1!��U�o�?ޯk�dXx"t��wA�dc9}�A�{�S����@>��*��tDS��b��<e�ɇ�H�]�}[b����8^��op=��4�= �?�9[�b�W��e@�7j�	_,1���K&�9�J�n>�.��<������Q�m
emIl�\7�%�x���f���m�r���͋�*�\��jsk�4������Ot�V5�1,�;��o��x`�-$�/�Ә�F�P��b�7���&�e�%�ŧ>F1�J��,:w�<�O3�� �y�1YQޛ�T������݃�=ѡ���h��f���m�
���M��Z��G�D�ǻ�|W:���{<e`�o��֬��5Y�Mi�/�pe�oc|}}a�N�{��
w9�͢~�+��D|lՄ�hq����G�3�����vsxh=yS�{:�#!��^����vB��E�(����9�R%�����J&��zeG�{�E4+v�Z����;�W�9�>dg�4�˿��9Y��q��l|�N��A�����O*�_��Ϫ�M�Ay���Ŏ��iQ�Į��JW͐2_��D{��{������M�T`f��C��[�S��(���|�Z�r_l,�`�e��53��#W��ROR-���[�Jl<J!���7wl�p�/�n�{5���(�^>����!ioNJD�餢`E���2�՟l�3TD�>Jf��Z�8�#�R��5�4�����0�����'���i�����_���)M�l)������!�j6nes��s=Z��+�3���ٗg�Y�IP�/�y��ce��q���si�������d��RQWN���nU��]�e����¦�����	�����	
[P0���L[�~��	z�����������%wFR�,��Fʍ���O�Άv;1�<A����!=�ۂ�R�I�V�/$�RM��0�Z��^��a��?s�T�K�I�VL�ӑƮ�lf�/B�->�l�/��O�'وN�S�O��Z�N�tS��@��rK�IԣV#fN�L}�$�Q�o��8���yO;]s{�cE�y�X���Rp���rM:���]�n٧f���kb�_�pS�<����j�P~�;e`�3�5�r���V�|/`zG����ϾA=7?�()Y���{��.���[��ݯ���Ӿͫ�I����ܠ�F*���Ƈ&n/�L������Y��Φ�Vz฿�˂����b�b���F9�0��}��5�������Q
c��R�%��E��=��/�t�[�Z��z&L�μ��,�m�ut�>��K�E�9u5=�2C��Ç������Ǆ����
����?d��"�)���o}�_������Zh�������������D>����o"���&��o"���&��o"���&��o"���Md�F����W���[���(s�ƫ��n��s֫l��>�� �rY'�����Đ�z?����IOl�����e���������V����_��&��o�	�&��o�	�&��o�	�*��������o�	�&��c�jW.G|��W'����v�v�&�@�����v
�%�K�(E_&����wyU��k�\m���������(ܾ��8�형�lL�����MtK���/��p���{����ȣ�ˮ��𳔓�/�Ô��WyC���`F*nn�_TT�O��z��EWp�g���
5��̢���G���#��8���Ƿ���7ӡ,��7�-�`�x�~��JB��׷ֽXu���p�C����*'�y˹m��jNӄ�@�Mo%j&7ה�_���[��"A����{�a݆��Ug)�����l��� �ɋ�|imfj�^�ݱ�ɉǺY��}#s��c�˨B����O�XK�Ǻ���U���6�-e��?^�&���h%��o��{QRRr#sS���u3.�k�5q\�Y<��ʲ�X��򔢬ۺ��Q���la~ў0��y�����\�Ù�}��e�w�<�j���gT���	�臢R{�FW�zH�����k~OϾ��w؝�[��X\r����A:䑳�w�)E	K[�>������3�ܧ<��}�@�E"�E��[�X�r���M�w#�Z��N����ػ��3,:� n�8F�f�LK0���$i�F�E9!�c(~�'�W��Kz�hg3�;A�s+k�!!h�ٯۈs�����ϫs���^�(��_7ISeŻi��گ����E՛�	3�.cJ�Xl�?]���DO�@
�9��Η'�eD�1�̾�(�b�������O1�)>-���\|~��(#���8����twKKKg�G�&�~4�\�H��m�Ǧ�{�ĸOHJ.f}Fˤ6��:H�?u��f��f�J��+!�O�����O~�Zز�6��HW,�ʚ2z�6�a��[�����&d���ę\����u R^�7���F���|���+�F����{�5^wY{3(NƁ���w#ΩUUUB�h�)�mX�R�M��_�˾D*4���>����rXU&.d�!(����ۜ%:k��)�*�*G-*C�5mڇ�/N����us̲p�������\]��G��'H]�h\��?e	{��җ\TUUW��AW#��]wumy�/%�t��)؂N-�NY �7w1R<�-�as���D��//�uY�L�Ѽ���T�f��Xu���ER�-w��/OY5M�y��`J��������n�Ͷ�3�e�D�d߂��r�5�S��U[UWW����}�e�y{����u�Dt�����3��Oi;1��%L�������^g�����(`E����`�؛7��m[����i�Y� �#q��Ν;o����A�,��&ƽjR��7�2qm�Z���R'qO�o�������gm� �<�������ϕ+�x0����Z$xq�D#yv95U$ ��[h�O`�WF��Ow�1��p��v��+�:�(�>k�ak�o�3v�8�lp�Ό�rqq�+`��􋰰p�9�.�9�ͷ���=O���n�ދ,z��{���CZ��Ζ����i�q��(+�۳���ʒ������G�1\*�cA'qϽ��=v�#D�T��l`�-{�i�����(����9�G�OJJ2�%�`�Nā�K�L��^���S�|���5�
ПgQU�YN3���}E�Q~ ��(m� 0�9�gb,��n�̒u��]\ḇ��;<&��&ɔm��b$�+J�� �^b�oꞚ��M� �	Fh��W�2'ǣ�#�/�q�)�.fx;��wqD�j�@�m%=� �̯�l�Ǭ]˲^���ƽ�T�VgM��~�yA��=afVzw�����(��e����A��S%y6����O�摈U߹�����D�k������OM��n`���j�U�B'�Kw�l�Nn�I_�x��Һ>H4�*��bۊ�"�2���6�@�:��$�+y7pI��`�k�vQ��.2Y�,�@	Ϸf�c ~9��ɝ�*����#(K"���>�\�돸hPL���C�y6	{P�v��+��ńF��Q�p4R����b�A俬6�/�N�k���A�#�L��VWW��X~0����)tҵ8������L`�L���@��������+�z��'�V/���U�� ﹐BٍT��U	���~A�H"�ވf՘�|i�/S	��0��[i���qUn�ḪaN"D�b�(�Z��"��Y䭱�,��=�� )W��4�.k㘪ś��I� ��x��/��ܹ�d�f\Ov�S��aPf�Å4d0g��Q������k��=�Î�Siii�ǿ�,���?��p�"��	�����}f�fà�,�:�=�o!�}*c��L�g���`���S�#)
�q���x�eӭp�"��}�36i	kU��q�0hmm��I��Z��&�y�0 �����)�����LY�(I6�	h���q�g���VlD�3ov.l� t���R�:�[�)��'Ѧ��"k������d��oġ�$�2b�¶i"�򼔔�s�t���]�Q�%�g]���\aQ|���e��I��&G��)M6���&?!�؋�<2�U����Xg����̩�Y�p�$�_tH�b�d�u��i��O�8*Y&x�T&L���}~077�m~eM��^'6%EGG���Z��kp��v;6�p8�cjΡ��&�R����=�m��:������+B�����!i/�y�J�s��Lp���Y�����d�yv�h'a."�Kn��)�ri� ���C}#�ə��P��xg";^
 W���/���򜄬R۸]v�DZ |g�j�Μ�8��̿tb�d�t�^�dG�Gi��
rHx�S��N���F�(��t��D=h�5n�]�R��S�����eP�g$N����B�2��^ߍq"�7��,yiF4,(����'�TE�n�F8`�ƅi%%�1{�T\�B��e&�z�S�&���ƛ����� m�Xޞ7>��~��.�Z)�62ȔA�2��od���Y29M�!�Ǚ�ϵ�N0|����ݛ%�w#*�ï6|����H��<v?j_!��,΋FN�_�Ci^x9&*���,��=6�*@��d��U�{Oq��ރG=�n����B���ߣ��ֲti�����i\��W���9�'!���n5K�Q@C	9I,�ȅF�}P)?���㛒zt�=t[��c�TY0��fxBL������ǲ,���z⦪��R���T�����ZSSS�g�Tg�X��g%A�蛙�Q'����mc�P�ؽ�Gi҇�1|>��S�$�wR�J(n<{琢��i���x�2V�^�N�,--�`"� ��+��v��+�A�Ӻ��u1�i�.�zK���5З=���� 4��Mi�� %���{OyA�sD<Sx���e�������kݠ�r@I^a�+4h�V����,7ۄ���j*��[����n�6H�g>�u��k�c���7�>��V��:��|/"�J�.2q�4���x��:;n��s��n�����>�|J��y�֌D�La.�"�'��R�	PǸe8�˝��!�
�7���<�H#	H�l�&
Q�vO|��C��6�.J��q�M�F���""͐�[��"���*�n����y�b�Ni�a?��d|3fX[#���&��F�}T\�#Җ�l$��<�j7���ꃲ'�J"����X�Ƣ9���������I�0��͵�Q���~S7V���2B[(W�Rm���m�"Ng�gC��<��]�`Z��v1O8�d�"k�Z��z�)=�PŮ��w� yh0ªk�gS��֎"`n�����y[�W�3W�͇�)M&��
0���~��,*;��Y������VDZ�\4�-�X|i��Y��r#�~++��$��@a.�Ir��|��r#[�!��{/T��N^��ld�h�}tɑ��7���/q(�����d�x\is0��6��)�K2J@7���ㄫs�LN��nwi��A{/������&&姱�I�^g^����%IԴHI��ӳ�ެ�PfB`=�.�27�,I&�������e���J@q�!�Ҟ��^�*6W���V!�@��-�jծ��(T[M���D�!�X�����m����Y��'0�D����g��FCM4��Q����ޗ�>'���ĺ>wo@�b�ߏ8���+b�M�q]��.��X-�٘4r7�f�	S?�b�-��yb)�s���j3�ld�S/<t� uU��)�%L�x�TD3��<�ǒ�Ⳮ��HW��O�L��.��=�ʍ�Q����§i ��LL|W���_#��<0��/��Ҥ�0 ����n��FEDA|�x���JT����u3��4�2&�����r��h�eh�M�z�%�dܹsg2 [�{��ø��J������+E�X�l�
	�(M���G���6hLU@�.\w���T��S�D�n�V��"KS*��q��W^0�8�F���������J:''��)ER�Z�V����fyJj�N�<<:a$�N�-���1K�3�o�`i�z�s�����m�����*}�6�]id\5>M |:�g�'WR�j���X��aZ�uO�Կ%�(����У��4�NBz�3��\; w�^����9���ݩ3O�\�8b���������%����;�t�@�e��2?>>�?Q'-
����U�8��$��˗�	�'1vbܫ$��$<�S����6�Gp_6��O)�+�gK��gH����0���;���c���&���R��OP:n�}�۵��'����kl�,��
O*v{*�F�\�6n`W����_� �w�2BQC^�������	l�T�x�΅��Ԓ��p0��fC�Ջ��3"�$`�̑Dq|���FǕ�����PR�T#����BZ�to�Q~Ď�dބ�4a�?:�2s ����6�B*Lbx~,N�ӕH��By��D�!�>�vۍ��ٗ�-7I#Ch��3JS��j�6�N�ҷng_����ݒ4�'&I;���ke��㠡&�� Ȃ�巐���@��/��07���F&`T��xc��}��d.,�qw� �Dժ��<����e�!�ۅq�Jh�ܐJ�򇩓�x}�+5e��7�6m�m(���&S�O�c9���8'���A���z/ GO���`!���\x��? ����sƨ�����D�?��W���8����d�Y�
����8��Q m�j��`ⵇh�nnn�K�������^�slhӗj��,�XIM�Xn�V�T��p��:����q���ڬ"����\vƟ�;J�҂���q�6:�y�������>���"���d�/�$J���W�V츭Z�B����Z��\�BT�e`�Mc����(-c>��ێ���I��7��o�\�^�+�ku�!�k{`rr�]|BBB
g�'�3��d�)3k�C���o`�8��J�y�����P�ո/c��_��@@E�L�F�U�/(+��5j�8�|AgK-� Y�4	��á����tn�����:y&�W��IQ��C���n�$��LC�6�+�}&���c���6H�cO@�yaÌ��\8���S�ƦqW���^K��'CCC���rK�_�Y����+=s�҄��<�Vttu'�;v`r3q��ϟ?71�����+��<��Kr
�j�%�s��C��Aǐ����y�$s��!������K	D�j�휩�-��(TX�:�U[�e�@���U�Fh��z�VE��{�@ ؏f�Ct�%[����?֑��A�>��+�(:2�����\��=IM�-�y)�Ҵ��s�$&6Vv7X� J~NR��o�"�2B�/�5�2%%��8�@��q��K���B~�\����%�6�?����b�%��i�0\����h�,������(-q`��o/�Ft?�Q�� yj�B��C[[{�0mN�u�V�f���&�V�[qs�?�z'�I>�m��ӟ0�\�Ч��KN��d�n�ֻ���㜜���$���w;�{�YFT����7���C7h����Nt	y0`�����U'�&o�cw�^Pwʓ)���k�͑�p�8�醟y��P����Cm���@C+]�z��Q���h��k0muK3� ��%���e|+�2����=�Η%%�M`��>a�Ά�m�-���3��@V�`��b���y� �%��2cz>jB��G�`��Aט_GG���R�ص�"���](�W���U�_60X)�4�A��/��f����%��Φ�[���\#%��}���4C��C�|�t;�zz�Z6��쮕f�$���.~<?������I\#�uy8d����h����e`���g^� �=�ow���z�о�y��U}}}:k�d�,� �[���鑰��E>�tL´�r�"�>��.�x���3Z$Q�ç��z�$��iw#.���D;QZ�Q���{腧�(��N���M�6�?ͻk(��ێ�O�C��~�� R��~
&`�*���DE˽mm'������(l|�w�V�$�&�bb����_�;<Y	0[m-)Bk�R0�����gձ���	�1ץ��+�� ����ˎ��z�GH�Gz ����.��\ns_��u��cD���k�-ΟQ=����e1��w�_��4���+���jN�&����n��ݿҷ���Ͽ�#�I�q��gǘ[�6J]��:���o����w��=־�䛜t��@�XI���ť�g�tn�5(\fb�%/��B�0O��0Vx�?CB\�#gv�e�0�(�\|h��VIՌ����(���<�}�����b����p�k��/�����qq~�87VXX��:���}���b���;��J� ��=>�������A��$U�ʇG���g9�ui@��wk�t�l�8D�w�����LΕ��ù�
�+�q�@��5��L Ns�@�$<�ʜ�9��{3U!"����%�e�_'п��1;J���i��Ũ��ַ��h�G���R^�J^�`n�(��.�`$���:=D(��S:�=Ϧ��l�*	B��M~�832*j�"ʚN���ƙ���YaU���2W_r�={��H���v�����I	�`Ȇ'�y�7L�͇����q��>���[�'�tpN�4&2��UN|�����D�Fg��f����5RM!R�A��٦g�f#K�Lvq�������K�ž�v�ymT�6c=�Sj��
�P�jhl,��`�FA��8��\��I���ir&�G�f\ll�����Rt�����4]��T1 �64�bk���qa2�9k�٣��4mR&:巉N�|En�����v����DvQQ�4�z��?����N�R�nL\7�.�u7$<\��ral�)}a����C�t�l��G(M�Q���b㔦�ؤ�V�I�b?�*v0i,P�8T�ґ+i�n?_[[G�#�~C	�P���V&P�vD�E�r"s��Wn��>*�r���K�?�Tys�뎹,�l��W}�Q����Ck��b����r��\_��vS�/�!͕�:=2��~�.���b@ ���N��7S}��=�MH(?¯�����P��EP\���n�5>m���Q���R�"(���x�-�f	�a��7<��c��t+|�$EVΪ�Rg�_�N-w�%hABټi��ߟ�(� m'X�Ej422*����C���eY"x�L�U�d"�8Y\�� jN4J��s(��:i�K�VM�I�Z�nr9/w��Zrs񔕼R �]l��R� �-W1P�ow|`ίk*�	�߅Y/��Tt%��?X�}x��xr+�E���H36:&�H$~�AP��e���yү$����Aۼr��=�h������@j���A��YZZb����� �j^�'�/A_R,�r�1,�.��/�!���� ObX\^/�(����@SX�.��	��ﱵA��\�y����6OT��p$�]��f,F@���lr���7#-۾��)��Հ/�0�ڃ(M� Y&G!�g������u�̍��Eg�9�Х������/^5l�;2q�|�t��,:�ejl���Q[2���9	��" x��;�'$%���L�m`Zy��]�u�K�C<...���U�|�#諹����C��?�X����j����62�}X(W�D��}Q��} ����CU�2�
�Eb�Џ�!y8Ya�@���t0VbC��X[��{J��
�Z�X?��y�6�J_�B���]	u's�t,kG��^J	r����2��2J
-c$�zJW((ӄbYId/�qU�j�w��ƺ
gE����I����ׇG���h�U�Do�FRDDĤ�����s��"E��_'+W� ,�� ���zʁ�`_��҅٪X#m��3[�0XWW��Jj�~WkHjjj�J%��e�9���޼�\��7:�6����V��K3�Wָ�J�\~f$␶���w�f(E$õ< ���D�o4�D�7���Ci�����ح�(ÂG}^|ޫ� ��&ps���U���g=]XX�3�7:�<���y3�G�*��U��+D�]���B���
@�%Q�W���ǰ�E�H�.[�/4�ɓ��Q��_���v��^����q?*�se�{�9Hr�nNN�������h��(���2�f5bi)����ӡ�:�-���=�:�'t��b�ER����&+)��4�w�<-�����J������4��6(	~�K�z'�0�xV�|��0��ߩy/�W��)����lx�-7�)��W�CNA����[�J^�M��z�7:A���{�� e$���"�	e"�U*�e�`/��Ao@y���R"��p�}�s���U���Z1�z�~����lC�ߘH���<q͞42�a%
���\���K�*ʃ��/��!Q�Y�6��H�����r�btt4��P#��b��Vu�	��>S����B���6b�|��E�n��V����ٶ5"�M��(ߓ���[+������J���� ѐ�ds�=�En���O�R����=N�M�j	���a��L�"��` ���3�l^���q[��В��~�Z* �߉�8�H��_+m"�R�6�@������ݒ("���H�&�-����@8��{=����{��0O�,�ۂ�KFAI�O.��#�}�y���t0�|�	��cz�}��z��Aj������bo�f	�c�}j�����ݹs�SO�gch �c{�E�to�DG$�*��K54j˯��@3�Y�L_�$ю�^�)��NC������%%�<����A<rj�-��p�P|	b�\�ٶ/K#8@��Y,��de��4*Uj�T�#����^�����sYд����͹�NL���3uĩ��<(ȏ��(�U�𮯡ۇ��%���f�T"��T��?[ZZ�ӟ?�B!���0��Y���@e~�����8Y�Zֳ�,355�s�
2�T�
�-�pY:Z�ϐ~��@�f@wg�v~^� h�<�Gg��K�e��T�8��y���S�L�E|!��v�~�2i-7�A�p��\�KLg�޽w�x-�ȟAЬ���i�B��"�J6��*�S����ZE���ǥVQQQ|�h%�R/��l��+55;X�K< ㋷�~���:&0�<��/�n��d�_�)(�-�J%)�1\H�V�l���MO�R`�����h!Y�������|#� �������^��JK�E�%���n�Y��f�A.Nd��!j��m�u?��g��� mHP�H���f�eA���i�[g���Ql��S��G�do9��\@J����뻻�>:1R`��7����R`��^Na$�F�/��X�����N#ᴸ'�LBw+�C*I�6f*��R>:����G��S�H ����������<k�^�nb�:����S�ՊW���Y��ô�u�ʴ��QJS ��KCf���$T	`h4�[?L�:w��T&������#�����
���fdNy���)W^�\�:x�H�'��Ǣ��B/��{�&Q�`���&�gym�5�~�'�z}����5�����p��O�����lT�^��ߓ���̿s��˷Z:�L��4"V�W�Ł~ о����UG�1؄T��S{����N��J�Ԫ�]��'�@酻*�؊q����?�'hO�,F)W��Zn���9=��4K����)��#YvL�0����V��%�C��y�g���ǝ��� �XE��suz!�]Q8�~=V"lh�mo�a>�$�� ��m[�hQޝ-����;��)�cǎ�I�v����p+!(<���P�>��i��n���s�N�V��pJ���.�$�@v)�"U�����!�1��?rf��5L4y��@Q�p�"n~l*\p�[iEx,z ?��<X"�\�;v�rp�f/�y�T��O{�����u��)+=|`�;u��H�9�E����ǈ��̋�6���1Gz������z���as��B1d.SWGgBj+��$+�?����T�������|;�R��[���˃��X����#}���u���W}��6O���5���3�C#r�����(E�Y�5��vpY�&i���OS�+R��w,������6��g�\��4�R��)��Ν;_����X�C�u���ʒǎ�N���S��a����@u0����P#�6�oB,�Qi�o�4 xu-�f�T�Q�hOQ��L��~#�ߞ�i����3,\����]-��&S}\Q�Ͻ܅Z���haG4�~HS����Y����f�eܜu�Im%i1�©���9�RiF #��ã�Ux��&���2�@�^�
�y{@T	�7C����>�#ӆ	���<l�z ����ܢ�9��N�[�'���=��R�8̿�Bf������(��
|�?9[�7J���j�T�3?;F&tnv�	h,�/�[��%��� q��;�;�<\#���QH�'N���36.3���Q����v�NUL+�t�:h�f�\���.S~�"��A�]�[��g6�FG`�#�'m@���}󺛑F^˺�����ss�Zr���U�c��@;]?YV���p�(/�X��� ��'�ɐɃ�*��9��@y�9���iu�Z'm���5< �٠0��a��@&jb���D��X��$��yo������1�s\E�2!
��~v>H1_��Mَ������rN'c�Ϲ���v��b� ����D6<hx�9�ďM�k�T������TL^�����|����ن�C��/{o���B3��
)|:�'������R(M�T�7,!�@�Dy�ܤ6�%�m:��\���,]��Q�;��z�|$�4Z�Sy��?��v刃�ٖa��i)NI�f�Q@��7���
Ӓ��x��)����~Z�j�:0�*��6Ee*�AAQqG�
deY�DA��j�4aɰ��(� K�,���w�r�������3�w��C_ov��1j����F�7���?4�J!E�
�^ǣCW����!�Ą�ҹR�/�k,8��o=G�[J��	��3����)�3}���}fUku��M_�p|\��=�%u,�c]Gkkk9�����AR�/ى��Q�MaRRXVRVfq_��n��Dg���anV:p#��w���e�M��Ōҋ\U�#z�\zh��Ǒ��=����g=���5P�l������	�g({�:�s�T_PA�Z��Bk����dp�����|wq!��Ǧ�#��5�?N�IS�8��0�Xy��{���\��s�[�g5�^⠅��6nV�jv�mX�(�x���\���#�������ǙuO@�WY���t�����e�n�f�� Eދ;>��K�y�C��� ��*'��s���P��E}�VnZ�5ZI��fY�s޻wo�@������}�?`:9ސ��t�޽�cy��I���?�s)��ܺt��/e����x��/\͝hD��9uy�����l��Ӟ�n{[���&SZ�s�����ㅀ��S�}6Z�!L��t`��t�vIFg4� , ��;��!@�:���r=2��xK��)3e#��i��ɂ�.�u|m1;;��4d䩅��+F����^3<6�������傕�5io��G���b�r(`�j	��Q��L�5Y���w���x��}�&¸t�̕���줾��] aT`p.=gc���vP�i�z�ܹ�{��>Ҳ0���Mj�ճ8��;ǜ={<�ѿ�����^h5'�ɚT�GsȀ�I��]�6U�Wj�����R�{wd/��<�@�G��g+�b6��*���o޼�B���V����" �X�y?źf�Kt+�f���>���т���w�)���K��#�u��8ٵ�<3Ea�.c4��[1d�|����U�cGM<�L��������n[mq���K�c�x�N��/h�=�I�P_�F*A����^�;d��f�MH��Iofһ��Z5?��3��_vLA�<�>{}u���%�θ�k�Wo����a�f%$h3�,�-Gx�P^���+D��#�^�w�Y��^*&"����TR�Ϳ$�n�u�3���P����F��K=�0��l���2:ԛ�M1�Ը��P���y ���0���֞�~<ߟǷ \�x�9C#������v�in%�?��ry<[�Zv�H�:2��?"���>Wa���qH������_��.![��٘0mu9}��]9��l^� � T�;a`�t+�t�l�B�s$��ߨq%�粓�<VR�vU���q6ױj�������[{��1שJ	�"H���1f�2�-�dXE�{C���	��򢷇��S�qZ0�ʺn��		
���:*� J�i]:`&�l���e�{W�1����?�]-\����Nj�Ff�C �*�`y0N�D�����nb]}L���hŀs�@*��:���߄�5}n%�v^��f�#j���B��}ł��ʲ]��1u����u/�&" �Kr"��Oѱ����<�=�fy��F��\�)����e��z���]Kv,�#��d_��`��
��,`�&J��8�߭�g�?��ӈ����B��^S}޿�j�,��$M�ka�S{���m�u�=�@�M�Z��4����)N[�\���F�%��}� �:��l���@�t�: ʤ��a�H��0��_��,܋aC6,X�[-�+��p�O�l�6�.<@�#me�IHxϭ�O���h��9@���ѐ��2Cn�Y����b�!gT;�P}��dY꽒�����.�~%�%i� u��TQ�~l[6�Y� ���GaŒ�{�����
�Gv�Q��mY�<���T�{)e�A����n���MK���nX\	��w���f�MZ��޽�4j���utܵ��/;��MG��Ka���>W�o��B?�ҭV_�.9����?M-޼��}�Ϝ��W[_�:k��)k���s+����By�[��۶�¬�?���l��fz� o���7|�����|Y��*nȻwʮ�׫�v��<~�5W�ox�CB�Z\i[[��D����|�f(��j�P�6��*Ca�&�*ԫ����ȍLG�l��4���[�y��־�	���/Ճ�c��|>�~d�s���J��X^dN�b��s���0!��P�HYc޼y��!j�� ����Q_f��QZ��]qs���ن�����f���Xu�ج�*⪪����^���d^s�ݳ�ɥ����2��6yp�nvke����'�����U�r�8�gb+�a���D]m����13739��:�8K��ϒ^7��.��9 ���5���#;�!���t���?����,omjXɴ����I���@-2�X�qʝ�� ś��k}����
�Z�^�\r��ms�^^jjW
�U'����Q�Za���ɸYI���U��s�����hů�~H�;H�������ޡ�pt4&�}C����+AS72�}.��B�ǭ�R
����c �^;PYӌ7U������DJ��F��G�k2�����ϐr�[f��t�1$�y&��>��S@�be�����ݟ�*S��:�fGj{5��Ǐc�mթ���&O�AH~(//_���#{�)璲�'��IN�[˘a����S��0���!��G�����|������] zl(+�ml���@sP�?�ĭV�?��ƄS���=��Fx���g���D_T����)L��r7��X��<i�-X��X���X� ��j���:��Xpa]�C��t#�����i�'���~yx�#\:�|}G��6��5�k�ɓ'W(#N'�n#B\�M����2m�z�ii�1E�el��~@"�0��������ξc��vWG(��Y���ř��7�%sY�Q��UX�?g�(��6�Uc���{ۈ��&�v,�u�%�����b"��&_/{482������3b��f&
F��\����w�%����P�����6>��%+�z~�,�$١Ƙ3g�z�	SXk�v��z�wO���8�"�Zq�~3�ʹ 2J��'��r�X�%w;-��P�6e+5����>���Tzk~�޽�0Ʋ�@iA���K�g҇����bw��\p��?�j��Q�d���+L�s|lǳ�m��}��R-s�[񈾩Dx���c}(���Gg='M���'�̭?e��(}��<�=ɷ�τ�z�|���=�Q�^gѓ��ȢR<�|r����~�X�Xga���6�N���U�X����V̍�b'cQ��]�w��1l���A>
W��+���1Vw)#�"&(��j���Ȍ<V1ŝ}��s7��S�l��u�SQQi��!�!W�^rH'��r�lʄ����l#TfLv�G[�Z����B�	ǽ��s~�����4�Y��d������&�j�n6	!�?�q�ܹ!1��8X�^�>q��! �2�kb��D<��0n`��V�6'�����O"4�w�q5�p��o�7V-���d��q^>��_��W����ɹ�/8���e)[g�k��q��]�x�bU%e����nL<چh����Y�s��m��|��3���s��5���`e_�� R]�(ɰ���5�����x�s��u�L|9j�m��k�ǭ��5"��^�Z��ו�V��E�h�/��>E5w��}/�5��. �B�j6�Eg��\���/WwՈ�))��Ʌ���?�Q>�E)+[��
cR��?>�zZ��n˱ts��0��F�r�X,�RS�YN�Jl-��G�=k���1���K�c?'W�:��yO��%�c���V|ށZ �1f�/N��x��8���L�q��3_(>y�孅&��3�u��SBe7�h�{�%y�������"tkx2N{d~(��sR��=G��ID�v�4�r�����lǗ昃\���Bz~L�:˖_���T���*'�[���$�C�����eDEJc郗�b�}��$���#�W<���k�XB� ����`�K����^�.����Q:���M�[�&�T�,�����~���U[o������Yqqq:'y����ku�	�2���=#�)z��l"!�"*�O`\oqnΪ�:�۸��Y�����@O�����+11��1�	4���B+ԧ�S��֬×Ń�f,��`#wvivY@(�F�c��z�/�xs:h&Ke�ps���$���e����>F���B)0Dq��atC����F�"K]YK\)I�j�Id�MW�l���7�*������_X�nxx�!"/��=��K���f��[��6l
�6�q���Jɷ8ڤ����o�Va�G�r+�r}��=�M���,�i����
��Ul����A ��l��Pl�g+4���9_ӁX�B�$v}�ZG9��Y5�hk���2��N�L�n~�=`�F����\J����e4�S3��9����D����8��4
R��֥\�������q�T@ů(&[�̖Bo��^�P�ۀA�O69�V�v6�]c�*1�"p��ڐQk�����%��hA<�}���E����L�h��@��0,꾥����+&��� ���u&L��$K�b�B'�%'"X
�oː��`<�!�T���W��u�A+�	B��<b]�d��VF�Az�e���-Jr���jʼ爪s�	��o�?oE���9�)?A��_�4v� �w�jߤH���c�X�q�\"�?�
:=$X�u�]���1���1�%�r��.{�H�-��w:�P�b�-�ލ7���/.���ת�M9�U��=gR�
1�cm�sZ��"?%T����D����rO,�(��,�z�h7����"	�MA%�����M�=����oH���t'MpZ�z��w=NH&��N�ژq���O�ѳ��ϯ��ɩ�O?��ƛ2x���^&#7QI�B_�4Xss��A/�@c�'M���c��5(��E4�*_����/����jb�:�7o���*6��5uZ�9߂�cʚ�X�y2�ܥd�GYǄ��i"�5c,�9zכ�_!_���[�Զ���?A��d����F��x�gr=��?�Q4)��.�V	����ty�)Z=e6��*=����V`�1��� ��)P�@�z�-��.ct=.��2�ɓ"Ui�7�ڤch�[
NOҘ���%���d�t����u��h�� -���b�#�wd��U��M�x��XA�ܓ�]��75�ɜ5셾�*��>��Fx��|B�ƂӪU�@n�k����h�Ն嘠:$AY,h����W�M(��C3���-	�ύ��'%'[̒������$>��*���x��@��퇥�qm�:�p�2�hy%R�[@�:��F�[c�J*P�ʔ�e��3������(!.dܘMO��f��h\�`9��4���	ǧ�������|�;D4D�.�st�����M���I�r�ZO��H��m�33�m��H1�ܸ��^�x0�[����J ��X5T����_�K�gүnuQku_�5����>W/�4b[���F�3�̝|��vE@]�qՍ7�7�=0)���e����c�*�t��<���^:jz����y�k��bo��W>����/w(79�S�C`ͤ�������56����������=!K�x���Z�w�o�L�~����P��hR<�i��Q��F|+,�믿b6�N rU��f�4E�c@D���P�R�]��L�	u�q��j�ف���ٳ�]8�d%�b��4;�wS���Q)ӡͯohwW��c�^��f�=��感sQ!�I���������������R6�������_Ϡ}�_�M_�1�Xԏ�o�ba{ �	z��(� �$)A��7[vlCK�7�����G�TVV~ĺn|�h?c��Z�sv�ЗN$�)*Z@+�.���*ӏ)8���;�<�y� 	o���@�6�O��>�%%3����&���ك�c����$�������U��
�FXJ#��r$����|�
_u�Q�Q1;9'+�ݝF��o�P���(�����2�|�U�'05��遁�J��P��照\\>��0�˳���U3���d(Gs�y�P�g� %Hq���$��Zn�\��!�!���v��Vj�`x�͟�4�n���d73V������i��j7`�h���.iZR� ��
���H�mA)B��u�g�r�= ���C5�i���,E˗->��k����Ѱ��'�bhG1�*٪��dܙ=�9�7m��E�?Kz�����N����cyFaaa���$���z%���  R�J�\���`1.A,E����飉�5d^��@�wQA�[����8=��ö�9�u9}Kq����p���f4� ϗ�� �|����y�UW�#Vg�&����;ȗH��5M���Eˇ�7�&?ߥ���%�8��PJO]�~���W�\H�-�2u���78��N4���fՊ����ki|��8GU׻�Q�0&R̎��X�0G1��C���.� ��JVp������9���pw|��9$y�7�-����|�X��`E=�8�"��>9��j0�,�Ӛ%��@>���A�Y��-%++�&��I��fn�,�A�A��rٓ�%�J2	��a5uS���Ji��h�Ϳ�d�� "��`]�xJ��2-7�ŉjkk�}�ҋޅu��N�ڙ��P����qf �#�����=������
]�N>ٶ䪡 ��W�&l�ީ��f�ٔ\�t���
;Ŗ��$��ݑ��}�gZ �i�D跋�s�U��s�Фxu��O��������\Z����{nC?]�ZO���Qs�i9�Gc7�'���$�L�#�����e�޲�S�g�}ǣr�@�rr�
zY�%�Z3��8dk�C��[��E>,WU��wb�~�N&�#^��o�u횗>kx+Z����޾�> b�kB)uL}�<��Ј���I�N�/�		�6��^x�;�#u��CG�{���3�-!�:�P�Q��|���P�������[(�*"�c$^G�1��q� ����Pw������?RRtv������Pr6F�\ �D�� �w�c��%=l�u��U�q|�YӰ*�^=J�>�%�h��}�@��)Q<x��C�����_s�2 ���s�|=MxLn4�s=}p���ӈ:�=rlI3�ʌn���Ŏ��M����I:Zo�|X����0+�ˉuOr�S�M�����z���t�!��.��.�����b?"�-�I��i��q��	�qTS�]���F,cw:�T�2��Q/tV�vq@#���V�
�5B���j-�7�ɚ���}C~3�����?O� |)���7Ѐ��{����y� �����/3`�{)~�A�儘2�y,O���r�${E��[W0h�U߁����x}v����g�(�n��&��\�`���jw��i@x݄�"�Z��cT��J��j.'�k�
�������Ƚ� '�}���<R��{�U?�u�@T��K�����(L�\�]�+�٬ex%��؈�Ox�4���s���,/���KӫG$��7�m<��Xڰ���8�P�����D�KG �۪S��D�ϡDI��%�y)ѹ����⌀���zW!��٭���z�XT	��!s�y�M��0�����\`���^U�A��5�-#~���0� ����y���K�q�oA��?��j� `���Q�J�@�A��1<7d
*Zt�2F�����c�d���ʠ�n
lNms��6'�UԚ:uj��;��d�{���G����_�q�e\�a0���-?d!��cµ�z���C�|=ߨ�k�o
bL�^��T��kwo8���rQ���_��0)��-���b[�BM.E=T�g��W2��!N�]�y�&�PF�'���	�yO�YQ����\�L��|����nj��f١�K�x��u�Q����ܔ P�����΄�� b��l��x8ڦ(L�tj��^j�����pQ�����=��#@���Y˅�n�d�vv�?0�G�J�y/=)1�b�2c~�m��k>�;bbߝi&E��?���Bk�(X������#���]�Q��u���߬G����sKp�{�ă�8D\��S�)����>V��f}�k+��-s��#PC?���c�#1�X�T^� Рq�r�<Iϗw�5���`��=�s���_�D�pM@�}�;�;����B�U��{�%��% \ރMixنl��"����֯c��B�7_���
-(�������C�$������X%b�!Sa���E��>�a?�I�"��th�jh�Z)>g����紧,Ƕ��(0��|I�ҙ�z��uV�7~s����nfZ]����3Sܸ�����=Z����1������;�K�҇����k#}răg�������]�0v�%�zI����X��&��X�&>��h��p=�t�0I|r��6yT�j� 9�R`�Đ�g�A�=��[O���gCX�9�ܖ��<0����r�z�:h�����X�x��%!���I�KC�Н��O����,�q{|�~�&;�i��g�+��\o���2|��j[�Pd*��$�$��80���?�
�ί�H�'���W2�Q��Z���>(��s&�p8�6C�&d�A[�45��CeZF�4�^���\���e��a!H!�4l�z"=-�A��$#��?�j�,S�`�|ve³��B�i-�����A,��3�M��o�mV� ���J��V�Q"�q��zL��������/I�������
]E:��[F/���!2a�ؑ�G_	����CPR��1��'�2 �7��H)D	�&����G_$��`�;�wX��? �6fP��L8���*����������G�����Hv�Ü$� �ig�62��{@��,��@�}����<�������[u-�R��Lg�����6�|��w٭-]�$���Jzc�,Z�7�'Bܛ0�Roo�� �\�`���8F/�6��MUn#GR=1�K |�8jc�����P8:�� 5��;�+�g��yCW�~.��18��XҚ�p����苮@�8�F(q�Y��BSz
��qC_����766����]V�����a&�Ka����"W@�qiii���}�OU�%W���聀���"# *hqޣ���kt'����a=�<�Q��u���~{|>w�Y�L�!��E=&œ�Nx��x����:^b�(�͕
�\���AZF��b�y1�i���cJR�qKvR��j���Zu�eh7R%h?����9/F�7V�+�8L��H+X,���J�u;��x�DQ�h�y̬��˝�ܴ@��;6L,� )_�״U	��4E�y}����gF�@����6	"��h˶R6W
��Φ=����eR���(kV}Ύ���zտ��hjz.c�^�M:��5�G��Ϡ��@͂"��_����6(NЧ�|[�~>=����,���J�~?�z�N~�	���)�͊���>º��ݤß�r�4J+��U�LE���Ķn��i�x@a��E�U��ڿ�rl����a̐e�F��iP*s���Z��ߨ-_�Y�č?]n�ә�I9��s- 7��ʊ+�_���K��9S�[(�?�I����5p��S�Xd�Y󯉵�_Y�ڀo�5�&qBޥ[Z�]�vt�a�ŭ��~Ox����b��åf0/�ا���p6��[�a|�� �Ԏ�XS�	�f-+!���dO���R$�m�[��:��XުG���*�J,�W=�!���A{g���]�-�K:6�F���Q�?���������c8�����Ol|�3�����!��3Q[��bd��
�Kp���Ƭ��Y��PK   ��{X A��?5 �J /   images/1a82a878-f7f8-4e20-9f5b-ecefcb5937dc.pngT{PU]�6��GZJA@ �(-"����tw�#*� ��-�twww�k��{g~fBX��k�����,>�}|y9��((�k((��`���>eT ����iأ��$B�P���R:H�;�Z;8���8;;�M����m���v&q;"�QP��K={��5�����L��n�z0I��}m"ii�����ExOx&��_�� ������hSO����
��(M7��ߣ�Q�H��=$�������[��ܹ�\%q��L���O<�c�Ċ����>G��@���s� �KG"3��	���^��
!��U���i�=�6o����E����D{��ܴw6��bݕ�2�a�����e�p`�p�/(\oz߽{p_XE�$�!`o�@��ȱ��HN�"�75�
�y}�ۃȍ]))��W>pzz��������dȦ8Ȍj��7C�����O���JVv�P�ob�N�I`0[v�5���Ϩ��ug!��k}��UI9��ddJ�spd���������}��-	)��۷�����8��\���R��5~���+[���$://�e<߹9��˳3�9:�q111L���e�L��Bu6���@�?777g����}B��Y���1�e���v�.�kS�$R..M[Jj�:���h�j�ʡ��ӈ/..���������*X��
��qAFJz=���q�+-�m��,'w��Ç�����������^�""�{{6 �kCّ��(,ял��n>�<h�!$��L_>�#-�J,�ƌ�a����V˟'p,����eQ\R������%Y�@>/((���%kddd.Z.y����QX�I��p�|���{���8%5�ȼW6JE;�� "�v#����:$��/�;$J��М�Z�>����橱����EF�^��Sn�6$��S?��fag�@C%%�~�$<<���F������3E��r���&�ֺ���W����Q9z���$BG����V�ҩS�P)��34|C>uy�k��9N����:��F�Ǳo��sqq�vt�C���ݸ[X����w�i�m�d-���T.���=K�>b�R�o���I$�)'K�������yyBo6<�����eB�+RG\H�'��I�Ҋo��w��2ڢ��I���%M-����Ã�;�X��v������̞dgg�m�d`d�RZ��u��O:?������۟�wn�%���ӝ�(cA]+�)��ÃKe�>Hdi4ԓ�o������p޹cхMBFVl>
��*/�oV}���w�G߶�/A�>�~�%ݟ(�>Y���d��K�^Q!��I��($�7?�r�B��辜���]�KKK�N[c�^�ᰰ��ed�IiMă��8�U�ƛ���C���5~(*]28���<G���I�?��
�u7��O�"�.��ہ�_Dd�����ί����I�Ʌy��؃ֺǛ��!��^Gøttt�����wqs�y�21�`�|�0��r���-E�h�%>V!3�-/��j������.O����2������֮��	__��~�T֟k�a�1��ۢ���^HV(�Z�D��Bس��?W���EK4�,--�5V��2���~T��b���W=wI@)��������_�	�Ll���5J�O�yF[A�۷�)S}P��PpK�u��D���0bE����+ Aع�t�������d���u��p��?11q�7*��i�<�@��� ��μ��P
�ܟngOL�Ia��נĎ�d���P`~�w�tu�q���\l�((���fy���b��%�s�O�ӄ) 9A;��;5M8�pO���@@_B���N�<c%�}��ξ<��0�xi1Q��t��}pp�b=[�NUI�K�/6����y�>oy1/�Lg?��J�meJ����e�˳��j�:���yO��K��ض�*3i��Q���p�/��ι�x�y�ssz�V�!]O���������8���+��¸��hw'D1-��=bb����T|�44�#~�/�~[�2�$꣰�B�&h���|���PO������
�=�����ǚ�>�<�d�22X��������GČ����,�������J�_����J��$1��Xv,����vT}E�`@��bi!9ϸ�Te�н�k!�::T�}_���hI8[����nJ1�a�s�9"&��\�$ l�W�]po����x�Xf5cb��i{B�����\�Õ޵�rd�T�N��`�M+�d�ޟ��zi�դ���p}�4�F}�*��9B�gk({�M�w47?1�׊���6����VE
f��\R�RąS�p>޾�!=}J���S`ўXa7/����b�=��e��ܷ!&F��B��^���5y��A62%�sC?B�>$�A`�r1�ƈ+	%	�}B�+��Eho�Jm}�x�(u�7+&ǫYg�Bv�/C����eH`�gg.2!�]��2O��W�b'}�d��PƶR��M���Wދ�o�v�����G�'RV�����bozzvY��|���c?���Pe�iU�s"�[t�j�d��%�Kk�P�F-��j��HII11/đ�j���Џ2��L1QQQ�hE�UV���prf�Lri �8{���XA,b��g��d���c'�
�,�V��^�i��<;+��T3�?<4X�����K�ɴG�E����#��y �T��X2�+�Ȼ�����o߼)t;6���`���6s�FywFiE®���g{�g��#e8�_��7��l5z(-5A%a��o"�5�J;��g�j5J�K�k�1W�*"��u=M$�J��`�����Hnj ����}@�P�]�S��2���$�r�w{_�!4M��Ǡ%�?.��[B���/�/q(ʉ��L۩�3��h�)���1�xGL&�iT.h�����M'���9����&����6 n۫c ��`�a�h���jm��D��O��$ٳ�Rur����n�і��V�2)<X�l��	#ײA�"ؑ�eI���C�ʀ��A�p9�FR���;j��j��`T�ڛv�Uy��N�@1�����K]]�斖�ؙi}��ů��W��77���c�M捷޾p\���:n�C���8<��Ch�ի-X���?%JX�ӌ �չ�������K��w.;�F�Ɔ�$ɓ/���w�ɗ�ҹ-I��[�p'%н��zC~��� ��Pts�6�*W�������;�����T�T�+�;��$�%YY�`z��W�UY�5�F� ���VJ�9!�B�l�Aݝg�#ɣ��w���\I ր�>��+����ݻ/��Wb�7�p����`v�?Y`M
�H�k��Kjs�~B�FF� ���&I11��;���S�=sp�bL3i�;:�^���椢���W=��j�N��Z1йJ?A'N��U��"^yjM�x4����λ:vvv�;���/���k�\8`����u��B6�� � �9'^�9-������;�4���.\`��6��u�'���e��P٫989� ���{�5$d�.|.��ݟ2�Q���F~��Yq,jd)%�ټ;˧�[��7
�[����PA{ׅ�âJ&�!��}���T������#���,��,�*���e4�ť�}�L�U���m��~��z�%�*�+1L�5`J�������R�;RQ���q�_}���b���$"�N乺��T�Ķʼh�,�ˍt^��}}+��b�-_�"��v/��_�U���+ F!��ǧ�9����ר�'>H�#�#�z���,|�߸Pe�88s�	����Ť+�8�{i@}��&��y?==�����g�O��	a��%�lA\�����5׭��6�4�|L�F��дp�[>zJ}��D�ځ��t�s�X����e�/6��id������Վ-���w�'ı3v��f=~mޓ�ҌD`�)7wK3~�I�%.��/vt*�� �A�9��i���2u6�~�
u6%�ћ/���mѬ��Y��^�tţ�G_U'\<$� ��B��~�ܗ@�����;Հ߭?��z�K�k܃�; �ߚ� ���Yp��� HJ��v��&5\o[�S����;�4-᳉`�U$"l@-�~w3X���G����ܭ�M�
��y�����M��Y�w�^���k&yᙍf+'��D*	e'Ý�`X�h�ZqJRBO�H⠛��gU0Ԙ�B:��̣0���T�(�P���%�n�_�-�8CCG/�xl�$���;Eߟx�G���2�_	B��Z_�Rǒלu#�a̂���v��z�/�@<Q��vs�P��4�m W��i: �]W8��j����l��-��ޝ'Cҭ�P(��Z�8cݾT��ެ=�0�QŜ�Db�nUT�:Kv��ӓı#�gP��H�����pCA��	�,���b,�������ܺ�YXx������۷���gD����̹G�n�WZJ�se׀�ߊ�ٳg��稾��8�L��'/�A��9])(Tn���%c��;��X��N2�=C]__W�I�	����|��K�d`�۵�CXj����fG��
�ly`�&`˝E���y8?�~�,K��zU�Bwo�i�e��+�~�j���4����A�-�w�ׇ�U%���8q�W>�(AԕjK�D�f�U�.�P�*�w(�i�Be�j�9�|��������򉀮X5M�jjd|q��� ͹>��P3f+�U^�Y����|��u�B�M�RjB �����Bnl_V�r���~�����6nZ0�1������W�^�!����+�������N�U�ߝ�ei��J��9XXvm��8��>��x�q����{O�+3�[�C�+ſ5�����<���M�2���������|\߾}���I��9~˃'O �����5�?~���_�+7��P��w�tr��$�{><������]�R��F�YL_(���b�i�o-.~JƦ��޺!�w��n��p}BCݽk;33���~��r|cs��zƣ�֖,�@�PP �p�	���R�̯����ԶY*��������n~�)��a��Dd)*��5ZFOaSs�蕌�NvY~b�H�	�nMל"SN?b``�����ӹ�2Yl����w�/r�G�y�yw[�UJ����6��R��E`4��GNA}u2�iz��;լM�
$u���I��<���.ZE�T%[�.�tJ�6
ڄӬ {�/p���C����)���9yy����#
,Q��V�^�	>;{��ˮ�L�����nxCP��M4P4�Q�\�>�O9��)tH�ީFU�E�J4T;�$,wGn�[ϊ�K��3�EE�8���ঝ���k�Ъ�������\\�ΰ��~�(6�e�(�([^ɣ��\��Gܜ�_��di$�TQ�|E�C.���@�͗�V�D�J�������^khh F��?=�1��X"�}{t�P\R���� h)YY�c�X�:7��@X)���6��Ɂ��@�WV�����h�����l��5�(��Q#O���*,L��0�W�^����N�[�Z�����"gNt��_�K����`�R*���1��=�I�RS�|�uM���u.�q	#�uOW��=\D"+�)) @��<�ag*�����|4�����W6R! ?�7�Z5�C�?���&��G\�$k`�)�463H\jeq��=>`�>�����\Z��y��`�u�')��k>* s/�wsppT;m���kkz�ř�~��]�Ls����U_���\ZZ��۷�������<hL��8<=]����� �{�!޿I�W�E&��27�ԺD9�V���w����ڣ�m'fm,{歈�h������UY�!���ya=U��k@ "�����m���_�n��|������3�����[�0Y��~�G�t��A��Y�ϟ�'��mܕ22b&ļ��8Aȑ��CT�V�v` �s@�[�z�O�ylL����.�Y'a���Y^���*���� h"�S=Nt��̡�77�C���̤)��RRS�?z���U��B��_-��5M�I-����P��]~YH�9~f����n|�mͻ�הL��ᯖ�>�/H � G�P���<�&���u=.{�Q����M[��(`3��>����V"R����<h�����w77,,؀��J7�� %҄I�i���n_���pP��@��]S|�*i,�~��-�f)2J�+�m�~����N�|+��G�ݻ7�$i���Y/����o�W���SW�qUW�T��u���襂ƕcU�?�����
3$Z����ao��*�~,�H��Pʹ�O]�!!��X}ro�f�ilZz��e�j'H������CiE��V�D{.���k������;˒�t�b��\��3Τ����h�HOo��뮮���A�JcQgP�;�~:1�w����g��������������O{�h�؎Հ��,%Ʒ1SD
R�>�ʳu�XM���\���^�L���"��֠����U��]΂�FV@����`yU���f�&��ρ9R��i����\z��~_�`ZF�Еb��D+��Vt/O��_��U1^�(�a�>?F#�Ł�2Z#�07g%��BC{λ��.�h�:��:��x� l�V��G ���=E���(�^8n�{":��X0<s�M3]>�5�s#Z��g�^^(�=x�S�*����=zg{����d+(���L���Pع����Ϊ����En�c����,&�;�Vq���������dd�q�|�=�_t]O���d	KH���(qY���ק���a}�-���	
��)��.�"�*��w �<�!���Dۡ�1����2�V'B��0��o&�l9�^�I,ʴ'C 4q�_��@/SS�^+c
,��>�����ߣ�;-+���R�3?z��Vԭ�P�v���[�
�I9q�nX�ږ�$� ��ժiIeyh�g=�S۱Rd�O{�0�oO��s�@O(�G�%%���枝���Z4x{���'���Ӳ}��$�/zJ}:�L���H0�DT�մ�g��ߍ�
�݄.y�7��Q��}��������j�ܕ��Y��˗ڋ�6��F#s,i���zOa##���}���z����ű��)~��n��b�A߷���`��Nн�{��<6G�98
V��c�)�\�Lqm477o�ޠ�Ry'X!��_��/h���7��%��~i��chP��#1 
M  �����eR���������i+f^��WWWƻ��9��Q���!�e��9v���*o�,����?Z��Tъp�D�RB���d�Vq���%[���YKe)-���
�F���n�edfvNɎ���}���s��,h���v���kp0#���%C����A�bCyI��� ��LJ��94����@�U_�k�R�q
4���^>6_��ȡT4��koa�s�=ƺ�Yr;��������J���$^�G'n��~�$�@2A��	����u�x���U���g�AD*���(ĽD��w�_(��F���e�6ܶ@?��`���ג~���J�vh��d���3[>k�?��?�N���B����b���^����a�&�%�>/���pC)�/���|eFz ���hE�T�5�-�]o��vjv�9�KL����3�$OON���	���<<=�Am���$�VL+.>�{���p��1[�f*�v1'9t�  �3����Y��	#�v�IJJ�l����]l���Q����ڕ�^�kc1_�,��H>?^�DRu��
��yYZ&Fƶ�ERRi�kD g�EH}��ѣ����<y�zR���i`���/�rs-�,��^_��oe��X �a<�&O-`Ә|C����%%%%>�Ƕ����	z	%��ĵ�)��L�:=<���;�&�UZ���Ǻ�<D	4�S�+"��X�����x񢳷W��'QPt���$\xe�ݻ�}ɒ���qg@���C��jמ	�����(�ߥكw��rݳ�x�	~�O_H-EC<ZM9k2�Ԕ�jDx�<T �����8��v*ώ����naY��cf��?����k2(lڒAw��Ng�Ł�p�V��FY���1^^Кi<�.5Ғ��lA���B\\H�i�ٗ�đ45����N4�n�M�w�OO3Anh�Z8�����)���{Ine�o�.�AG�ԣ���3��7�-G���ׯ_Gz��C@�2��lt�5���r����*�i����?��J<(��C	����!L�{?^(��3=λT���݂[����p����(�t)A���5�i5U��3��b�6�+���vQl���p@����c��Fu��o��/8~sE���]�����k�G�lBd����ņ���P^^^1F��������v< v��������|�)��rU���v��+?���u����-���F�������8��c3%�e$3W�T��3�N��r�N2k�y�8�:��fT�7@!�q4�fT}�j$��*�Π��z��]#\qI+��r!#���t�#{udF�������f�U�:�#�ֽ�������XC��8�4B���")�:)��Ss�s�ݙ�㵵��V�/JqU�և�(tqLLL�Y��;�ӥ�i��*iO�*嘃�u��'n�RE���J��=�˄K__ML���
KJ8���p����p�g=%�[Sfdll�r�dҺbM����Ç"<݀P�jqq�~�P�U�uֆ_$5����\P��4��;k���V�x�?�HP^���0ؾ�����C��M�~H���:���~���m?n���j$_[��*_�t|�	h�����Qr��l�d��H���x���4[��&�~���p�p2�t�is�#7��jͨ����<oo��xv�MN�����ݲ����kP�!��pŕ��G� g��I���y�KHR�����
jhhxoB�5]զ@=��w�Y;E<��]_ko�
LS_�6�4#xӒ�Y"�a��:�kG�$ ���ޞ�PUQ��������x4Fĵ7�J���E} ����ED�++ ?Ň�p��s:m�gL����9	Rha{�g|��2���`��*��M�7�;&�?ح��ɜ�����В�`��3x�=9�}tvW�Sf� �� z&&,�T�t������K�3���>�
�;S�:��(^U�r���;�4$���@W9�beP`�ŭ�~������-j�W����4W���=wp����ݝsN� ����T�r��c�|����z��(��rE��g���e����`���*�����Ɋ���\�K�������A%�^��)f~�(YZ���:.�9�)��0���O�X
ׇ����6����Y�+�+[�9����7�~���,xV���F�d;�9/j��|-���edDDE�6 xR�Uo캕b���VO��Zj����m����-�N�����@�{�e��䊉-���3"H��7YTLth&C|�]�0q]V�M�!�/e^1�vvOA/�<�%$\F�po�	�b�ks$Ϡ=��(UP �#s�w�o���3ewȮ͙|���"�e�Nȸ�5���t]ިo����t���T ��@-���5e�PX���C���$��aÉq[ ����Div۩��?1����>�K��k�k�]L
-B6;�0B@�i��N;s���'+�*�Ip�<�u6��4$�ߝ�4c����F ��+1`G� B��?�M����8[="'&n18�]l%VΝ��9�7�D�#�H�Ҳ�׮�V�gy`�
ϖ ���U�������(�Q+�����S��o�Sb~�yx|����
��J�*�y��`SW3�I]��Z�?M[���˕���1;�rxU���;�*�H$�͛7Pm�W������ j��. M�Õ���դ���Z�S'P�@W̯���9���5�Ƹ�*���m������)� ]�H�§?w�z;[J��=��Ix�"���gC-�;+ف뫫�9_�ʣ�o=���.:��Q]D�\���x� D�ľmLo���ܝi[�G�U8����dR��YQ!�t���V��
1�c"����� P�^��8�Ò� �k/wj�(�������<�~_۔�� ؋�ѣV���N��w���UK��Ltz�X?[���D@�t�?�ks��&g����H�I��J;$7H�ze��(��~�H�L��ue�@��AEG��\�30|u^g����0�n�d�]�no�(L�-7�xU����� B��in��c	��؄mc
,e�c�L%G���F%�.���U (��gb���n'[�%��b熉.Ww�ě|t�4�nʺ?!+�G�������=a�E�_��j�Ut���C�������ɓfc��|�����?��S��8$vuw>�Ų�������;4�Ԕ���#�����&_���x��.����*�|q�d3���mvs�de0l��ѓ{i����UoE��Π�������Oh��<�P���'�V4z����+�QX67���>d_,Ο���6 ,K0)�t�S�I��+�V�(������o3+{�[�
ܱm'~���Է�:�_l�,f=Oi@�\�+#�T��G������ڗp��A7MC�+��N��m�EG��4�+9��L��$�	�=�k�P�����4��j䨒��9���8k*�a߿�}�VU/3�~���\N�<+���b%^d-����Z�}- �R�1���RS#���ߥ�����,���4P�xtb񍍍+��2�G)��i4@&l�ŏ�%��6�<�6��i�@��3�JI���Yߦ�߻�l��n���L����!s,�#(�����
}��.{~��[�����mЋ�������ֈ9�D0{0	�p�?����'̙ix`��[e�XTT�w��Sz}��L�ߌ�3��'܂���{dd+�c ���9��	�j�_?W|�y�����Z4�)�'.W����&�z�2oZ��<���'��������Q Ŋ��h�Mck���G�	�3.���VX����?���'�<��h�^�����"�槂;Qh�jcv~zzzO�5�a�l"�չ���8��X�tS�b��##�Ք�������r�@W<jkOg3��o��5v����wxp�́�`��flU�8R7K5��А����*�ͫӝiP���Ϟ�"λuՋ>|	|]��yyb��;��{���aҟ(
�1ٞ(S��	?::��E���^S5x�D�4��.��U���&SdD��aR
!YgddԲi�9���Vv~����`}qqq�p�Έ�Hmʹ��L���\݆z+{�^1b���5��XN��z|6gA���񮡽-�%U\��O\�y䕔2~�<7�Z�]��J"7r�q<���0�L�_>���L�����(P/��m�t�MKlS��;y>r�@*Y�3Y���=�蹣1�J��~�CY���6� ��i~�N�iI;���j6����>n��޽�3u��5����JK#�D�����1�hݗY� R��:R9��<�����x#����+�h�/����|��~ �7u�dekhO;mk�	��;�޹�S9I��b���|��i���sӬw�3�>ѓ?�yk>]����bbb�lWi����"@T��o�Ԋ�O�^((�l����I���ߞ���:��z�cF�z	���p�r�bH���tׯ��ɨ�$����Z(i�vq��S[6��zXJ�U�\�����/d��) ��������nf��]<t���b��`��T�I)^��۷����ᜨ��Yi�����?ֳս�6�¦t})M9�j�j�h64�[CeEťD��W ���D2�"�����c�Q4��[i��U_>�ʮUf���[#X�OD� �Ur�2
�N ��
���*﩯pҳ���)�ɧȠ噘��::;�ͤ1	���JxK�'##���̤b����%%���j�*f��Vb�WQ�<�K֥����Ԅ7��c������>��,�痏�W��*�D�i_�������zy݄M��V+��֞����]3��xԍ����As���%&���W����ִ�<����7e�k𫆳��Oqpp�ܽk;�3me����^��g��f5JGSP�:����!q���s��E���{���bk�+P����� |�AdeJjj�!1O�p@O(ɍ�YLW����<��P����[wm��{b7;q�����$�g�BO���D{�	ʷ|�eĳ��*Z�ݸb���g	P�,�*��@�fAC��`��T���1,�+��K,'��/ded"����Ѡ�g�t1�&��\�<�$$n��2,�냞��$ 8g����8��"ԁhCtl�����W![�۽o�i��XO���SHY�����E��b}0�H�%����J�CG���=ҵ���z��꓅ֳb�	����S�,J9x�����]�̥�?���@�=/���qZ�9ԕ޸�?
��=��{����J䲧���c�rƻI��7S m+v�=0�Ų�22~yo]�}��ڃ�㔅�C\+�n{��A6��qsM�y�ߡ��>^Z]gcڙ���@��'�s~a���g#�AD�:zg�.�����d9��	O�t��;l�ҳ��D}l���8�\ܹ�Gbb���7v%����w�+6{�����`��o�8D�\c��C�z�mԳh6�3�{��U�;5�.8��p?�<���b�2MO�v������/�V���	aAG��_Z%����<(ILN���tu}�ϼ� �զǳW2���{j�ZQ]h�"�/��߅��C[z��懑�~ɸ�G��@�%��-8�]D��̷w������~����!n�6��l�ʠ�����^�M"��҄�����z�i� �4".N�ؘ	��W/��@ژǪ�"ʚ���i;�~����?��vn������I��f�~_�~���k]�I� >�~r���zohP�渝�:��@��+

䰙�_����C����O�^�w�������#�T44� nm�"2L_��˙���Ĺ��
�Ǚ����͈Żmd���4.Sla:�T~����֪u��mX#	"L�KK��0ME�����.-���s�@��5��̌�l��t@�̂���7333Gk[��Ch���3(d,#�6�̹f�k	���¹m]j�F^5�U�>R�o
� �>}�����Ľ=�z�.j*��?e��^{:�N0��	^�����*�ľ��&�z�{�՗L�,���۩���>y�l�o诟>�������?N���`�pߟqߵ�f��|����L��"��CZ�2���t��|5_�������Ӿ]���6���w�Bb�2���?ɒ��y7&+�3p��VOv����5���$�� %�M����W����zrW@K"�y\���3�ԅ�,�1�=M���*Ӭr^��>��y՚]Y\�������)) 	�Y����K�wrb|�1ܛ�c�����!/''7}���DT4�F��H���{�(xj��ɦښI	���ڗ��,wc�&�̧c^@{b ���`s�Q�ӝ^�0	jn�I�����@��#r;�x���-���#���*::ؒ+.w�ɫ�����O"N+#}��^��uX�}�͑���]]]4n#� z㕶����**0�J~����ƌ���
g�hj^��6���G�>���q0e�rJl�S���Р܉���!E��+$!���� ܵ�������@�Y�����\5���0�Rw�~�U��e8^������=A��x^Sc.Ŕ�$�$=۪V&`�;=�P&�^����܋է���,j�����A��2^�Qo�KZX��V��v��=���.��w��������pqq��G޿���y��ɯ���O�O�d
�����a��Ƿ��r

-������xo�\X�w*�WtX�J��& �A����K�v�����!;�祓sT��.MMM�!�#�@N�8��&g:�BEE�IO:?\%&"�cqlgx|�Ԗ՞������Gw/��rNLae�e���5Ԣ¡z6��@M�m�C��	�Rбq�`[�kǀ-����B蹸¹���_����IL��t��w�"v	�]E6Q`ۉ2���bT+8��I���pH��%''��N�U~����?.�k�CI�B�k�>��)�K2R��o߆�:���d'����7���WL$�7������Bv���lzigqs����5ަ�.\qy(�ʕX���N�����'e�$�����+Y&�j��:;<G�wtdV���Ƴh�PC�,5��,�G����k( ���q� h��¹9=�9v�xV��ufrF3*���b=3.�YGKK�ήx�/d�ڑ�b�k2|5-��X D������D11�:#%�S�`�Z�ܑH�O���r����E�������tMnd����-�$%6�7--�R�N]���F��-{�S<N�h4��R�5)0ۡ��:���&�O��A:5}BC	Eݎ>+���1��M�[���S���
�~uu԰��V�5y0��㩶z��z���)�W��4mj.��w��feO��ס���B�6�����+���O���XЃ!�u`p�VV��; U���Y�Cc��v�E�Ĭ�Y�����!P������b�x� ��.���_�z�	$%�\26�_�����Q��w�.���4���^b�@O�����.�F�L�7��k�95P\�߼}˵Y���Y����_�3=�$�wzj]��Ԡ#�hc([I�yn^�R�������R��SMPTթSy;P���Mn��ԉ�ŏ_1��4I������@��蚒]-�8����e#�����<̾s��DsıoG ��¹lr�۷o��M2���""�����	��O���#:���Ui�X����UTC�ￄ���+m�� �t�L���/")i�"�8H��=I?|*-���{n��&&����/d.�>�ࣂȫ��*..����e$�� V�u����#ҵ׺hL�>c~�:���3-�_��	=���nnn���v�ﮣC{�����1bbK�ʼ�M��߿��A��i�'G3����Ŗ��D�I�;ZM���l�!}Ϣ�S85��r,��RC]��;��qq�AɸEZZ�%_�«������r���Tvvv".����/O��	Mdkd�
&@�V�i�dP�.�L�K��6>w�m��B7B�2'�<�A@������|*������gc�M]]~`��%b@~q[���-�)�^��z���
���qӀ102�(��(J9��5N�׳����P�a��x��f����(�P<�lV��v?9$Z�ޅ�r��L�����ULnC�W�lz%�K�ǳ>�Ꭶ/|&�/^w�@p�4W�NU0D�iǡ�{ ��@@�Ji�����/ �BAA�t�>N�)�am�AP/-e|RRhR�n	Îl�UE������j@"��(x�z�v�D��tvp�i��1a}�u�8���qEw�ڗhX\��"�'@S���|3���;�����&�Hm�0Y������b�|b�m�L�����0�~��S٧�;	��v&����+l�a���W�V�[*�C$���S���S�P~��~��粧������1$��_Y:���?���ά[>�,��C�,$$��	Ǡf;y�0�'v���i�ť�H���_���^J98�T��=i:�1 f陮H�qɼ6���U�`����������ql0��%�~4��I�b�w����Г�y�����Q3+��A+����"!!�<r[�FE���8����NL�T��z��Vݽ{W����r�ׯ_s��P�����Hݡ��ө��AF|4� *�*�]z���z{�S;uh�C�	Uۀ8:��M��%aX����	4?��]+���ۢ7�K�Pl��u�x�-(�΍H�?ռ�����{O�Qx�p˾�� 3X���I�XDDD|�t�;�!p�)`�n=N����+A�&����ˀ��1��h�[���js�dV6QSJ�O�P��T��&Zi(�j�b�+�v��_d5-���^*��40����x�P�)��͡�i���4+��<�H�s�?awo\oVv�3 �y�w�.`���kor�fd&{��:�ϑE�GI��.���(O�hJL�W����P۽H�;:�Y�W&;/D(���ɵ���e���=}�&�9£fe)�~� S�I�G��7��g��h��ju��ϛES�F�@Pd�����~����X!*��Q2�$����{��![[���*���~���O(b�_�����G��k� i�������+��r5�f��<U	5Dx�G�:�aw�ʞ9�k�8?�ť��3���G���Ņ�n��m�m��|p�s������ÎeeeD�цX	(-,>�b��?�������>驄I�9�^P��ՙm�0����LP  $�k�������SG��e�q�&��X^��&�cckV�o]qq[zBM虙3SU[^ͻ��!=p��O�H�{v����ʄ6�p��RBϓ`,�YYr'rNJJ���%ffm��NZ��g*%�	���hhh�1+�~���_�q�������v���i�Gs��/�aa��˫��J���<4��C�񐃃�_�?XCz=;�F�S�%�>.6��lO��+��`��b�m�ʊ�{
��*I�NJ�������Z��ӎ7�������n�5����s�qA�BL��d�+������@�ۮ�5�[��3�Ξ� %]P9N��%a�Ąx�1V���QǏ�o}�A�Yʤ��"�rH���d/�r"��|��o�!%4j\�P\|6�`?a��_J:��g��(�����|��u��?�w�&!B��s�z�oѤ��'�5�~P��N��<R�$���Im
���t{�n�Py�j���b��a! ��|/�"�C�N��2�-�D{Ⱥ*@�W�����͎���[9Ðo�&���٣UjA;���X@,�}
?���l�m!}��Sf>�RV����ޞ{csFJ�\������zڱ9Z����m	u�1w�V@��<��I�t*��0翉nC���qi9o� 	�S1��I�<�w�|�JRE%|�
�n��ߟ�2;K��wD�22�pΈ�	EP��(�k"�p�	P�SQq�=����+ǟ��Sۇ�xb22?��/�kΧ�*::!»�ē��B�r��YY!UG���8�ޟ��'kz�81Gi]Q\�g��"b���mwU���'�`G�C�D��A�,w>=�,*���Vd�Aԃx���\�u}C�ȂC~]sM&�)	���j�c�V��Vaqͬ���٠�.נ�ż��fP۵��ƹ�ޞ��ָ����4&��4�I�c�����ִХ�qBa�r�ݎP:Y#�t��:`)=M~�St�"Z	�{���TM��G��Ĩ���x��$/�W�>Ч���KsŔn�.��D�6�j�:�����؎�x-��m���5X�~(K����0���s:��7׫�O2���FF���q��QU5�ߗ�F@�AEBJ$	i)�K���)�n����4�����z׺�@�L���=s��� 7'L��WO�<���937w��xo�ӄ�N�,]�s��$DA�U(Rp4�+%���0WK�&�޸q�j��^�
���u���CN4��$�Oê�U'^1�#���7g�� KK��Ȩ8�;<�å��p�!7:>�v�X�����M�{�&|��]޷��9?wP��"�]�����0���l�P T����%�{��1F	D&!-�G����ӛ߭��� (�Sa���e�@iu�y������� !̿q��v�?*�NZ�����#I��_/�6�׸�W�7� !�T��45S���`=�D�8(֦�0a4�����ȀjG��XVV�S�U�_����Ә�&J�i���..����{ KMΎv��-se��~pQ`���0�_��$`Sb�8$�6�s�|q~�Us�
�V;�*z�z����E�'�h����Kߩ{����}K{�f��fKB��&��������l@R�wd��_~����r ���IAo<�g2�����ii`�W����p��kR�س�>��� <z��C���=C���=R22��5X8;7��X��%l���v����D$N��r ���k��ދ��|��h��[�S�}��d	�w����ɑ�Q����g��ŧ�1t�&vN�a�r�=����9",w�{ �MV_%��ƾ��WD\�-Y�y���y�cv%;I��*qY�������@{	(0�$�zc��2ʶ/:C3���3�ÃZGo���q"6߅Y��HFM�[e5:�;≁�1\`���'�s�����3�2jO���r���G��U[[[k[[>���+zԋ��,�D�V9�Vz��,�^�~%×2P��6z' �(BLC����b%�Ұ�h�eWQ�C9�>`��$���v[�L�ܰ��JN7���[ṫ�������w�Y�o�0^	c����~+�bM�#QQڜ�.�ck�0��?~�<h����@���Q2	�Oj������z�H��B�D������'zލ��ڛ�����(�{os�z!qOd�r�ʚ777h�bM�C5��=�r}�I2�t��k���)�h<���J*bN�C��-����?���8~�D�}�ݯP�  UL���$�W�o�U���6�il�o�}�f�B��0X @���x?�L���eJ@���K� V_�ش�SV��,�U�3�(f���_^<�*�n�ѷ���k�<]"*=���XJ�(��M�&� lXf^^�,����ŵ}��~v����[��N�����y����Ui��p31�dee�Kp��a�Sp�X��kaR`�ѣJO_#t����+yW0�Mx3Ktb"A��]���R*@�w	��3A�,���ר�P�&�QYIK@@`/���{�/��u�~aCӃ��$*ݾ�(g&�K��O7�x0���<5���?�2���e8�E�{��H�6=��1Q�ٳ��bԗ�ǋ4\���H��_��(n#*�($w6"�O���-u&���WS�jem]ߓ��xAK��uy����5 +����C�Z��II��J��{,ym��V�_"q䱏��p����^!�*�ʢ%�"]���u����ijɒ@��u&�O�'Wy�@ ��q� ��X��z�dRW�%�ܬ �NV0�e!8��LF� ����f�u�7�1���Afgg�[)TLm=k�BN��*�U��,��+r�����ư��yFV{p��E��M�����Jj�����6tpd��&�|�3�u�wA�����s�SP�%w
�(~O#�H��NP�����ʃ�>M
W���/t^������ ���/��a�������N[K���Dх� \��)wp�H�w�o�ՅM�b�f�������� ϼ����߿�t���7,v���I�����i��W��� �CF����>j0 ~�7Iplg��	�_�
pw{ip� ����3!�O*�s�
�QcT3d�����Z��ŧ�
		������NI��d!Jy���&z��T���w���V�����\�%PI�6"��ܧ�*R*��<.n��d��D�K ��K�Eb�x�� hR���i�����\؝��e�m�&{UnY�^����
nn��q���R�C4���d�ɋ��hg��x1^���'f�<����X~Jt����U�l^8�]���F_ϭY4�M��A��7�����{�,�>QW�Y�M�Cꀵ���E��ԋ���̼��.w�����"�B��O��F�Lq��Q�B!��aa2a��4ef.�{n�O�.59^7�R�7Q>L+�WA ��������o�7�[b5h�ٔ��v�7A{,|�� ��C�I���ɃF�Cuu��U-�xP��'����Od��!��'6±�/|�6Y�/p��Óp]�m�w�xm���AsAsU�3��c!P��޽kH~%U��1ќ��S��͗r��դ΋�W����("��H��r��Z��x�U��v�H%�`)�����>|_I';]��]�ء3Q�rm(iq�]r�2���i������vS�t�k�@��x�)Rh󽳹�%��,-37�|O@�����zka���κ�TZ䜞Q3�I�r�xzzz�Χ��w�7x����p�i��r�l��|i�Ke�Z}�&�S7�h)E�P����O��[�Ptw�]Վ���6�p8����]���~NG �MQQ2��\.󔆆F0��V	vvL��u��΁Ǚ c�}v�8��y�홸glX�}���l�4����&xwE��8*.��>�u,3㨫�+=|����r�YA���aj�A� ��d�Y���<�u�@��M����}W��X�j+�{�����sg�O���m&_���7.�5�Ӻs떌��T��`�{���s��MIޠݡ!v�f�&�-�ˆ�`�� ��m�a��֍�.z'�OG�0#����iY"��1�W2��L��Kvv9��h�F�m>�=5����SE~�`*@��=K��揢"��|S�r�Rt��p2���􍛇�}��ΪWp�,C[ɸ�
��L��k��N�G���*775�۷o���o�8�'O�D�^�y�9�֢O���C�ۈH��1�������Z�џ?ߊwM���V�<�
�qnv^5��Q���҇�Sss;Y��;:�r1�1�n� \�h���'�'�6�YZY��"�BcbHyB�
N��?~�x��	�X���p/�n��%��j�U��~S��)57tTn����Y�H��$�pK�N��~qcSS[���N̺zz7�Z�+��\���@IƸpQ��$���������,�T�ax���+Q):jR�0!�� �J=�鯘=�ݗ/@��� �`�C��:U#�]5�XFu����~�N��6l��MX�a��[���@��e����ۈ�h���#�,���]֖��t��a���FN��[^G3�;mɭ�@MC�eǺ����ΪQ�f�T��
���0Wr�Pk��H{^��瘝ʼ���H�&�/����%��uX��>$j<yo�=,h��0)ޒ�����=��L����F"����o6���8�j*���\A{�:9�x��rr)��� �p�B�Mn�����m��e�9W�n�%t*�0W0d�J��2[Ԁx;���k�4��@�t��y�)y8�㴴��{������%�9�5#ƅ#�^�8iG��F�*z�moӞ4��>qW"��-��Qn�N=t�P@P�U���nG�����n��ט%�n��L\����kpXsY�#1�oO	�Ys��7dG�-�oC�~qNg=���ʪ�X�Т�)/�;6�bgb�۷�m"i��RR����g˲	➽/�*QG6B����;I��Y��N���N�_�$.�!�Pq��C�Ž������� ^t�Yp�gQ8L/)*���m�ρ*��ˈ�Of+���/��g����G{�ө�X�=@��[�0c���j�;az�����w[�0�5Z�顀D�	����
�nD�}�=��b��h�����E�E��������j0����E*O��@Lس: �f9�򃟭�J\��e����ļ0�p=<,�͔�?�_�$%��� }�P`����{��|�	r�%���<�*�����'�vvw%�vM���K�-��V�qf4��I�Ύ梨���mY];���*�g�}j1RQ���,<<D>19�12uqXR��CG��dMf������(h�9Ď8,�J�X7�G+���/&=��]��aZߊ�gmm��s�L-Q0&A��C�]1����#�bQ830d�d�_a��(�  U�N�A��������=��W�}HH���9���j�ƺ�UJ%��w����@'�$��쇶��'Ч%A[���<�̄h�(0sss*�)G����5o߹#�������ɰb���T������P�!�H�S={�t9-|��oJj갮O��:�5��'��|<8�2��kW�!<e�2YHIIͶ�K����3��.�,f�$eut��i�� M�Y�Z�3��%�4��p}7H& ��H���s�h�b���f2;�<��.|�6"BƮ"���p$jt4�� ׈HGGtVkM���\���d�1j@���@@��/�T>�0e��hҐ>�$Q�/N�!�^�TWӳ�_	����|����o�ȿ��U���"�[�wE2��n��h��L|f�D�lVΩZ�ؽ?2��[�@��w�آL�.�U��ʢl`��;0:�
�4��D�N��U�u����/�L'���0�k�����8�%7�.ȉ��<�-�Η* f� %6��\Ej��_�x�+Eƫ��_�U�>F���pvq!���+�H.��4��ڣ�+��h���W�eH�KI�z�c�ט�|�S����}���֋m��D�)cGV��(�_�K�E������X6rpPK��ዩ6��b,��Jw�G�ba���7����-Q�V��.�fVF�y��$Ǳ�S���{��P^.
���������ˮ�HB�K"i�XJ|i�n�7X��ZƫbU�� \v[R�^!]ݹ�����tl
�\M�~�2d)̗>|���������L܄7���L�bӠ�X�MYY�}������	�l0#v�*�Mp�1��g��w�<|�]�	m2�2m�;�]� t�G0�%�	C�����f�j����s���I��������M,"z�g�>@����ٓ����O�i�����~��FGG�;�
��N�#�q�{Yı۾�G^o�g�ϛ�ڶ���T%�z���o����d�������ӧ���VW�w�F�U��Q}kBŇwz Zш1`��hl�5b�_��� Q~\࢕� � q�F%�s_�t�������o���?z�h���@�0��*�ti�}�U7��.333�����{ T���u������'�w��~�"���I4��.��)�r^������JBC1���x��Y����\o�恅�uQ�	�M�uq��G�S�� G� � ��Fх�8@���Bn��q��m]bJ�] ��wމv��x������������%�����O�.�f�y��Wv=�������W]!�י��Ѩb�n�>@a�#�φ��p ��~Lt㪱����t��xk;�4v�WzK+��]�q�!�}�Yt��:= ��\�탆<�\IP�~���,v�8_K�~�����<�k�G�&�&�c�����ѫO�>��I��	��?8}��B��D��/���n3p- ?��(X[�XO�4}�G��!�V!}>!�:��� �oQ�� o�� ��cN�Fq���R,�i� �x=���4�gϞ)E���̴0��ii}��M9v6��]"CTQQ�jN��Z��1.+;�hE�tm�/hZc�����j��ȗ��v��~K/A���Y�y�~����7m��)Ⲩ�1��`gפ��??<�Uk�H�݅�DOH�5J&�h����&�U/o��h����1*u���Mz��msB��8�u;w���*�*���w#iEz{�f�a$�=�A�R(	�;��K���Ŧ��iTz��޳Cu�!qy���� A�b��(��[���풑o"��b�@�\��mY�i:��pc,�eIաY�������q��X>��o��kiQXt&��HMM�:gV#��I���&�O��G�F���^u	Q)C���:�|�y
w�ԫ��Ք!u��]p��kn���.T�G�C��Ru1)��=��'kѱ�KWM��?x���G52T�J������V�����|)g''��*`gm�������V�_��Ȕ�`�ta�t��D�/81�� �(�W��ʑc�B⻭,��J�*��h<���u�"��7��I�E�}fc?89$�A�"ݧ����)����ѣ�+z� �di�@���vyq�3j��֙���܏Eǡ��8Zl#&���Q�!0$<F ��Cޗ��<Xו��}L����g�{���B�wՠw�x=��GD���~����N��s��,�tW�����\5��EOOO�KsMhA�=ІT�q]F����-r
��J���G��b�2ԲD�"1܃�g�.�������|��#��	��p�LKCeQ�\ﯚ�cgbBqY���idd�;����s��F��k���~G��_,���y�x��ۣ�F	��'G�	hx�m��ɾƯ;ڙ3_�N	�
U����@W�	s4�E�wzP��:kB�K��k�����s~r��aaafp���� 2��[��
F_�㝎b�Sec\�:�Ǐ�^��t
�����h�)�,���~h��]`:���Q�o
��2t�F���B���%�A�{K��=J�Y99�G(�ξW�tZ�Ɵ��c�����P�\���	~�6X��c5��fff�ՊU��P��ӟ�����ثc����GfN��2�N�����5`��U|��6@̻@g�����]BEw`��9?E��
V��nv���YFn��״$9�I]���+�rpU���\+4�G��
JJ�y2�Ń��{@�AW;d>�Zn߀���v��3mm�+"��¶��0c�*$�B��<����aĆv��Ց@aA�
@Ã^VyK-��yܢ0��r�[1X�|�Җ\�9�-�_?JÇ���Sr�����F��]���v�D� &�v����O�0 ��V���5�gZZ���9Zs�_�渗k�#i�'��n��h��v�+=*SC��&ҭ%�&r-�Xn��P3���c*~���v�B��xD��o���a?�m=�M�EVGR�P$�0��48(\�2�41z�愰��+�IY�J���}��*�w�oU�U������2XJ��ލ��#\�̪|�6���!�K�K��Ĵܓ�����O_���d�4��E92��♦fY����$zZr�`��w�H�p��6�`E7���el`�:�p�-�G M�=v�8Xz����Gi=�P�/è��Ĥ�~����w���_�P������7["�4�$�?�`cg�LW��D�`e%cg��l"�d��G::�MFߕ���K��ϑ=��Aj�����I9 �\,:��@^�<��J	PG�A�ehSW�aigW,��k�
��'��]8&u]й���f�;||$ }\��ji���T�ګ���˃�֕m4��L�! ݢ�u�uW��!s�IBM��:��%�x=�+++W:�C5�X~*N�g�.,,p�	�����@�a/�L��%�P�Fi�s��V]?J�V��%`�d���!���]�>d O���Լ�E�l�(�Km�wl�����9��c�1�1S�<_�o�t���˼�+�}À02���BzBFK<qD ^�����h9�	�ǅ*� ��SRj��-�w>��,F@@��
��	U�h�\���]�r���NUW��6&�T^s8���'l���ҟnzr�*+jV��N��}U��7���'_��ls���j;$���K�0���".%�iv��Ed��_!	���G���,[rc,�<N��K����[&���&N@>7�a��ʝIQ�#���Цן#����ȯ�"����y�[�񰉈Zң9�
	����,H>?{cZ(0VA�{d����C
�Yh�󿌕�`�uN�X�M��}��K����E`m���o6.\|J1~�m��N�}p��$��Q�f-Э�!�;<ϟ?�u͜�ps+��X*����e0;,�]�0�����ǔ�*EXʆ}��ڠ'?��H�a� k�����Th�qK�=�$#W_�Т��i��Y�Z��V2L�������_7�}�U���b���A�5[��˂��2��Â��%���]�.��H��jV���p�������L`�1��v#��R��'U������e?�{y����1P�Ơ��:*<w]8�.�m��#�<���<kA�����\-����N��/�uE�r�$�364ƿ�G��/�C�bb�o�ٖ|���{F.!�b*	��y�g�|��o� p3�e6�Pv#�����Lc�:T���7�/���>x4��,�Q����\���u��˰���%ӭ�*::�|�V_IiXI�F�'��W-���b�����f4y�/���"낱�#�55�L�K+'3ʒE��Q�W�qw���=Rk��ȡۯ,�g� ]FZ_?a�h�:&z�r��pbL��	>~�ȝWl�����+�ڈ�s�l��[",�qN.�>s];�M	OC yq�*��vAa!��',
�j�-`� �Q}�dॺ9 #��/�bѮ�
����������O%L���mgppPub��z඀�p����C�)�H�۳��Z�����d;Z�����5�����|�Oqy�(t��������-B�1��_@����Hx������k"nC=�p��C{w�|���;������y7>>
���l�Yh�M���Y f��>��{||<Ծb(g�G�#Ցl��4�����K�k6��D^��&|m}��yyy�����?�\0aW�R��x�r��!O{{{>P\��@?�B:	��|&+=�`̽���/�����u�́���ϟ�LK�l�q)(�W�?����_�T���S����.\�9)h�ި��ڹ��;�t0/�ɳ�8'��"�1a��%�JZ«��557? Fos�|��3�Umm�44޷����v.�a֦�c�܅f�������5o��wn�%;�f�\��oR? `jɒc%@�Q�1���MFk�%��S�J�A��6㼟?�)d;���EB�(�hڼ?�;�<�>fk�
y7��5k�:��HN�{����z%YU��Q�ԣ�[!H�T��N�������%����wR�̚-��z��O��!޼��ִK�M_,�N��o�\�q5�"?���&�'ߦXR�9��O*�WO]�0z��d��/�����p�#n��aܼ��?5���Ve��]�L��<��ۈ��t/��_�� @l�h�d>SL9�g�̗|�,�u�v:)�O/N��D��TCG1�ա��.G$�痂%��w�VX 45>���seyy���m�'\�'�XK2��)b�I�i�׃pt�8y{���ms�[)C矅M��mG�����|���JI��M��K�3�k)���D~�$T�w�{�����v�6��%wW�R:�43��xX��h�h�a:�M^<��B�wvn�����,�����#&Nw����ѳ�xmP�z�uڰu�űl��T�{z�ZZ:�O�����P��~���D�d�8��qEU�+�+��S\�伥�tJB���6�(/����z΂ǹ�>����9�)��n� �Ûc��R�b��`[��Bo�����	��99���i�V6���OV�A0�py��ƧN����ʮ.�������b(QY|E��l�i﹵����S�����6�2���Z4"^�� �T��^��e��{�@*Ԇ{��Ӡ|����ޫc=�������0���_~\�y)`]XDGG� ����P>�ڮ��Zd�b[�I����'�Z߄�)v%I�/�l�a��'����$ �����~G3�{[rH���l�$Ď�U������]�� ] �3��i2^�8JB�	ҭt)ɛ����Z���e���B�X=��z8'���R��כ6�?�ݻ��c�ڢ���3��u�*ڟJ�>a>�3,��gϜ�ȲP�Ҋ���:1 �$�<D����{%s��v�9 7\��tb�����K�f�Mn�q�~~��Y�=L�$p����˷`~�?�����5c)��6-���8��?���ԏ��l<���������X)��hk̠�X�M��'�ڙ���?��R	�C����
��8����g��aQ?X��X�H�SIJ���v�O��*����oZ��11�bKeKI�NN�`9�KK�_��4��H�&������U`h4g�\:u���*`���n�mE�M��/yb`���������<�P[.��~.C�ũ��NV>�i!�f��� i�5��О�4����k'<�������r���5�1�mf��#��d��,�@R����E]��]7�*z���QMXޕ�
T����|kt������U�ɉ�f(.���=�*i��K�o����y���))>f��Q�l(To�����E�R�/�sPFQ�ZX|�mYh�Რ��&��zϿ���b:� ����V*�G����}�f�Ο?�i˽��Bv\\\C�Yo���8X��[�x}ݍeZ��C3��W�f,Wm���cJ�!((ȝ�7>��n췛+6]|���,�s\�����<��k����r�0��f��,�� 8*6+�T[Z�#᫪�..��0�5g����M��sJ�����X9�begt�u�����(��2S�H�܍?������Iq�a(�1�)�Ӝ��k��f��z��H��£+��3l%�.�j��8S�H�Д��ˏX�k0����\�F�^s�u15���{Q�g̖���5'7���D�"��9>Ԟs�Dr��0�,��©�om*�^�ȯ^�~�5Z��ˣ��<�V8�S��{.��OZCC�%��&�"9����]���bלC�����H)��/.\���͚K�u⇑�ŸS��TӑPAJ^���w��c�%�[���|��)F��%�� �	�˭،����}�a�b���<�s��|����E��Ye���[X�`9�G4G��gO��W�C���D�3�X�T�����i���s�s">%�N����� ��ʊ�z�\�jb}�U����Ǐ?���ee��7Fz�ܷ���*�ިTf���Y4�� I���9�'C��3*u����z��nƺr{���ld�#��aÌG~�����O̝c������;ڼ��&�@� ���3��X�B �[����ͦ��)b��[c%�)ʉC�"�X�����_�ʁ᫩�bP��l��
�����TMMz:MT\;�m~��]r����F���@$�c��/�����U�%,KP�w�����ڂ�����kۆ���͛+����S���%a1�_�8�[��,Q�8�oM�O��{�͢�ڟe�=�_O��-�Ȗ~�m�ɫ����Ύ)�Zi�� �|ϊ([k{�ڲc��D��+���ï��@�-e
Rd�<�Z&��W�^3�S������wF��{A���Q��vv��X�=;���pn��_]]�ׅ.��#@	FQ�DYf�ȠDw$��6;����s]˔��۪�{ٵ�R����M��������?���c�B�\:vZ�?�tr�t���Z�=^�����y�'Рn2��>|x��������_F�GGB��NNN�������l�,,���v�Bo�%F'ߢ8�l$��-G�O�N��t�./�%��=b�@9Z+;D5/4���=� {@�M#�D�c��h���(\#�B㎮��k��3���$$�X��(���-�쪦��0����ҁ��U\�p�QR%Y�<h�����nN���4pP9Yiю
��K2�.'J����Í1��p�A�����ةq$���1��m2^�^_�1�4�b/0�q,%�>�N�[{�[�U�6���B�{<����7�T63㨨�O~Dpf�1�r�X7�������W0bE�1��5��Q*pX��䀌�8�sF]x@��ϟ@<�=��ba �Mb��uv�@�Z{�.�_hh^,�x237!�����߾-���"�������~�z�- ���u� h��~�1	�S��zO����3����H&�Q��{H��<�Ú�-U;����i[�����{"X�ĺ��8*�o�ry�"J]�|�X�X�Sv�O�%v}�����$��Y��-��@AP�7�P/%�RNϬ���|�o���<'KDo�xM�H�.sz��1A����F+(M�Ȉ��M�]qt	�{z���y�`��|[S4�s,��׸8�W�^)E.-.�N�NӃ ���P^]���>Akk��s�����5���I�w�+�@���-�����Ո\F1���������RN߄���ޘ��{��eb ��SNX����p�z�k�˓�����PB�X�T�x�e{�D�{��X���c�� У+��s�"aJM�	�I<��c�ǎy��޻��&�DD�,���'��y�iK$th�9��֢/����l'�-h�5��S�3�������2
���'Y�7�B��ژ�;�[��yyi�����z\�� �eԘ��=j�w�*�ᦤO�X�8�	����@�$)wc��\:<�d��@�$MK�5��c/V��D�;d�&��ƞ��N��k�1-v!'�8oK�;S���8 ���O �dk�����<��t3�s�t�fk�XI_�A��
{i��ـ��O��ߴXD�(V>WE�E!�{�\��u�(�_��BL(�9�c�@RF|����W8��j���'�#�,9v���o�v��\�R(���p}�� dPR��
q���u�Fvv�l��媅uE�S~k���~��lU����eK*| �D\S23� )��n�@�/��)��N��{�˔�`��{ M������Ċ��Dt�M4����.t�33J+�&��In��m�ɑ�˼�����q�Q�4��������d .6[L����1�A���[�Y	d3T�J����`�S/�Z*�h<N�`��6�����8K�U99Jb22���o�?�L+*z�a���5f\�E���p~z:�4�Z���s�������Rut��H}/2���1�����J���1y+�:���t�`s��[n_Ns'*h��`'�4����z�@��ٮ�Ӟh�����wi�i�?u
�� ���~�$#ADD��f���\N�����XA��� � h�~V�4�gp�K�P�A_���7a�U�K�=o~>X�B��r�=�68�$����*������ Q�u�(K�Fߤ����H��P��޺3$-���;���Vf"QB/>BYEZI'�DV�ՀuH�YЈ������츻vF�i؈�k�G��#��=�����<���X@�~�x����b��D��y� |����ݪ��F9r
�?Z�Dr��n-�O�ZZ�,͇�M���a&F=�Q��Ӓ=M�`��9m3cВ8�8j��5�֙E�Nw���O�EEE)߲n޽�aie8:l�~r��eֳۖE���#�������n�]��U:I���b�3O�i�9�K"LI��������O�>u����P3�����򫬏�Զ�`�3�E1R߱���A��j�%�t	�Zi��W�q$�+���i�@q y\l�]�[A����1A�=��$�P��'�� ��� g*�FMM�����E�i��-o����Ѱׯ_�u���b�	�[
0�<O~�Nb-uv���R�NS�vW����\5��$=���W�h��ZA�>Nt�ʲ��j�A��DL��>u��qW�R�s��p���J�q��-������H�]�Y,(�����]s�1;��G��ܟ�cب��I"���ޔ�_죆�2�f�������#GW�����)�h%?��a��b Ƥ�9��h6)h�J���0''(��U?:�lMV�o�O2�bb{|��)}��ZZ?9}`��
���쨰]wNn���)?�H@���d�)ݛ+�9�,m-����y��b9f�{�b˕fjJLJ�����տz�5�x�;z
9�߹-)����^��S�{�pӫJѝ�U>�������������%��2(M��E����'E�ǽ�n�����Bo�Z���wb�V��I�LO�Y�=ݺI�������:�2��e��pk��*8x����w{S	)�е������ņٚ����1���lL[���䐩��uv匾r�__��8�ki`�/�8��.�<�A�> �[��ds�p��_S���#+��Fԕ����*���7RR��~��㆒��"Y_�_�$�R�Ô�����b-��<Oj���$ N?�{Tl3���\��i���A�2}�R���s���W�Ga����۸S.�M϶u��z{I����ت��M�Gb����;�0�1���!Zf3?�����;�p���Z��'�W�/�	�Yz�l��>��a����7~a��RA�@�PQ��Φ-ʶ��׌h��|��{w���?��P��nP�g#eX����aق:1���׳�NH{��J��JS��}.yu�&�al���{�d2��Ď�8E2��
�ք�e��4-��F��{���,�H��#�'�A��y��b��5}��gl{y��3�&h�F��Whh��Oc{��)������ӷa��5=eq���<9�0)BA���VXP�~x>��1a}U�M5N��L.�Ւ�qK�]o2��H��Z���I��0ݵ����mpڸ6}|��.c̨�ݍE�� ��{��܂l?v4d�_�����Ř��>A�EIs�؂�M<���H�o���"ai�BRQ�g��<'XX|��c[�V������]].�b$n��]����?-��z"'�|���@a�1s�E�FN�c܆m3~`��H�l���:8<�j?�z��|Ú
Oa��V����j�fI����Tu���\�-�l�H��ڨ�^2�r���:||"�O�U�����(�ai�w����h�yyO�>��$���}I�dvFY����\���b9�~⊆��*�����g���h��ι,��D��\HT��l\\r:�S>گ�������ni�X@���s����\*���靈"���7��2�����^���eo��+S�Ħ(�lda����1�#yh�!����[o�������E��ڒկ�t~�=��{n؜_�#��OBd��$`b�q{�=h�K��\�������������9�}���*�V8'{0/��UP���%'9Rɦ{�
W�Z��Eu�l挵���kI&�{#�f�j����|b[-�Jw��>�~��R��<���D_���17u2X�R������%}vIE����T�k���)yR8 �K�ִȘK�h��h,,�H$J��}�"��h��P.Kl��"�oOq��[��2��T7��*�\��G1���n�/�>���m�|�q��x��)2k��Ny�S�X���+0����|����ʝ]���?�V)��^}^�J���7��Z�G�����<��x?�S���|�f�H2]"�cv��;��R!�{栘a��{��)4֧�I����{/��������������p�7:��{c��o�n�H���1��@�4����;Z�x	�.(.Jd@s�Q���`4nB+O�l�v
֥Ʃ�g�<�:�����מ	S�i��\_8KY��jY�ψ
�P�~]������ ��TL�4z�i��CCX��=ϲ�έ[���ӂa����g�İ�=K��c��d2���ؘ�C�.n0�����^���p������P�,`���?
�ք0ܷ���2���}fk=�����|o��L��y�m3I��?r���b�n�K_mY����Nz��̣r1� A���lV/�d�KV9�D53��q[����1s&���>��[��N"i-�$��@ȭnm�v!�/���r����Gi�����jˍb���y�-%�*׸��E���r��v�^�ME{1�."�5�¹���Ɠ�,ySQ3U���F�� ~��qd$ǵ���&r�k&��P}D��P�(��&��Ӛ��`������MVk�qEF���z����)��Y��_���};��Q�����ٽcΏ5"s��8�K�-��09̎�)�F?�	�u\:qafF�ʨ!�A˛r�sL�-�5s���z�����?�6'�#��R�q}qV�m	~��QUήun'%[�[���|Y1.>�'���M�1� �	�I<c��);V����u�bp��$$n��?�	�c�t}����i��/.�˽�~�Y<�R�Mq��_��\˴J��b�c�����>�-�9�#�k���J���6�0��{���뙔��Ta�@j������)�P��l�Oo)=�iiuVs�~���qG���M�t�"�=���{�Q�@��$��ΘؾDo�H����د��VO�o컊Fdu4�7!��f�嬁?ǜ��w�ݢ/=Y��8�F��'���g�t^�c�~�W�<��+������/-�y�'y �D�~��	�>���"s�
а����D����=��s�bt��(�U�n�q���@ɐ���e�+��n���S�c.����w�M���w2|�_�v �K�}��g�C 1���k[ݲ����+u^y���'Z؅�rw:��I�3��W�-Ό
2u�w�7�����:�wfB��e؉�0�<,2�ijw����.zG��LH�$^�A ́��-�dN�Ӭ�Έx H������^ָCRU�G��!�=�J�,�^o��yyD1� �+jN���z0������Vګ:�x�I��177����������OY^��|����75^)1�eO��]6�R�S3����R>�rE��XD+n�*GP]��rқ�5)��������홺`,��ϻ�����"���R�GT8��.�~����C�E�|�L�0����e�q�5BC㾒E/�ؕ}�q�z'�!�C��tb��ܚ��ȿ�1��č��b��(xG!/��a���ڧU��?�[��: ٕ��u���lƟ�l�A����|$�w��/O��Ξ�q��Y�9��],�r�+^��a�z���Y���ڒݚ��h�d�]_R�S��@��	%BA{ق���iY�r���^��N��h����t,����Om��.�䞧p>rc� ���,0�Dv�1�^mzrc��D�����(��N���K�CB|*ɱ@�%���״��`�e��ڣo1 ��eo/#����cB�����#��������*耠b��o絺�N�2B�|�+9�~\`�	(.Kl�#991և�^n������ �e@�����wS.�'Bx����<����d�v��.�uQ�v��xU�|�h��8��A�@�ݥY<A0x�K�+sA&�Ɖ�C��?�*�Ԧ��)[_ês#e�>(�s9s0���\m��c/�1� �+v�h�܏qocv<�%FKEE�hg.`��x���vX9�{�>��0��5���~$پ$l�/��U�@c�		�ftm��*7��x�*Ĩҽ�ڈ�����������y� % ��*%KJ��t,H#��ݍ4�����Ңt
K������,�!%�﬿���'��ى��cΜs��AûY�=���YB�N�5�Z�EbaÇ� M7C.�����#���mK雸]u�@zw��V~9�� ��o�/{gO�"�zW����^Z����7�_�K;�1n�f�f��D��]R3��@��9��ݻ/��6]��*�ni �޽u�k0�1/�${�w��8�t���> X��#�J��i ��,�텨Պ@֏�SqK4�r��jP@�l��O�|���#x��Q���Q���-���ɖ~���}�K����qi��B]V�l�a'�oΘ�3����BW���]�Y�"��
n9s��}��ܟ��B\CV��B/>#�?�޲jdϷ��
��w� �G'1�ð�up�y���ڸ����c�R��YB��W]b`pi���D�&Z]m�[��ꐼ��9Ց�
��ҁ�ӯ� K�o�C�œT�1sC�p��u�ط �byyű�H�w^3׽mv�_���gN�(��P�
m��/
�
����2,��H:�4Y-R虨q�b��6ה������B ʘ�'�����ː)4����. 0���� -;�������F
%� ��z��zM��H�����u� �iǓy]EE�.i�y̫��Ю/K�߭��(z�5}�/����L
:��\F(��q��c�G�Y'I���d
�ʾ)J*�ꖖ�����1���l��9��q����݂i ���-�D�����B���/�6�N��`�!����ct��55��g��|��e�%�Fv�����<��?!�ۂ�
7çX�̤_�H�EcĄ]��R�����a����g]DV^m���UjM�>ҟ�+���	��h��l��^������n�M�]L�+��lr��3�1�TCh��b��v�-ʟ�`%���U�������>2-�%��I�m�c6qg�̞�L�^f{���C}R:��˻5�k8�-�(��:��/�8�<j�a 93tN�V��;Qt�yrر�E�W���`S������O�շ&49�þ��޾�" ���8���i�n[��c�E
��u�K./yT̀?
["��C���Fv ||�'��xQ��~ݝ^y&%
�t��ƞ;�<�^2���ޭ;5j�'���v�VW���gY�}n�PF��vod$>�+�޽����� -3� �h��LŇ��G�	d�*d�;л�vz���ptB{ƞ��ux�H�\Kb��B�;�}鬣���#�	���oK���p�eכc�<�Hѱ<��De��7�aQ�^�lU���D�U*�/#�l�ߠn;�s��?������C 	���da��_#4�"7?���G��v��VXw�+�s��=&�s|��4ٻm5�y��=z���u���������K�7�+Ӧ�?$�Rw�X#Xi($!���p2��G� ��]Ad���&��s�2sXut� ��L��_�K�Uq���܇5�{�|�����V�M!g������Ғ(���(8�<�\��blU��Z2�@�'�x�b�篳��������n���0+)4�\�`1n�3뛛�į5n5�^MS6	8�4��J�<��K2�B��g��j�0=^�V%W�̔����H�DBO���޿����^prz�&�oR�91|k5���yUg墤���4H]F���D+D1�aA��]��{	�_��)V�!�0��3�[vT��"Q'08�@&���4Ĭ�`�ƫ�6(wr;�6r�ӄ{zf���uѡ�Ɠ%��$*;E�Z�jC�� V��\�Z��r�<\������[)/���Z��ʳB	��+��OHm�t5౭=��3��7������LgnÛ������觰-�8)�FCJ�����(u�ھ�����8�:sscX6�I�re�`:ܪ �^�&~��J��.֢Q�\�t'�d�4_&/S��u�%�/��7�~���4��K����H<3W�jO��\�(�:ױ�Ʒ�$�������d�.uQ?#w`��y�n�C�3%R�W�6�t"��}\# ݑ�w�n�gkH��>�f�P�$��j���%�|�(Ҭ�,����ܡ�i�H�4X6�omc�0Xgs=��e
M�N����dR���+$��Ҳ�f^hG� ��|ʞNN9H�ܵp�4y���y5
~=ɣ�?</p�`Z'P�<z�(���if���(h�w��H�#��1�a�U"m�p2�������g>��m�'"{�8YhƦ��ct�$;���������+��'�T�Ro�+*͟k��Z��Q�21���_Q�r�\,x4��d�>�������eV�!f�#�rq�Ə^����<�WpmT�,;KeNnLfr'��j��6���}��oL���U>��O��!�l�e��?��ޏ�d#G_ѷ:A2�7�uTh������K�w�Q{0R_qYߣ��Rc���������7`'��goF���&ߥ���a��]Z��,���>,�N\i���D�9Y����W��@��	�-̙,�2����~'h%9�aV�N����R7�5��$$+%�V8�
�?������J�����>Lȯ�z��0����Ͷ����k�7h-f�Z���޸�d2ƻ�𫣇�"'t*�G�N���*����Ç,�ͤC�C ��Ӹ�}�z���BB�:��#�
�w��[~)�@4k�p�+~*���e��ަ>%3��B�lm�D^��dd Pl�IY����.��)x��2K'�.��MTy��Z���01a��|�"�E����F>�1c��.)�W����,k���$eW�MPBoB�D긞����n(��=���@�l���!�^AC#n��yq����о}��5��ڎɅ�L�Ь��!�k��?Z��R����(���:������Qj?N�D���9At^8�%=F�sSq���ig��ˎʑ
�����Xʻ~��F����/���A��fG�G�\����~T�N�� �r]���TZ��5%�ғ�k�����,͠�:󏽡���B'�1H�t��"UZW��M�k�Y�#�D�Q�;�(���d1�Y�i�{��ܳ��	������I���'�J�%Þ�"�d��̊K�K���4�(��k��b�\x	��)֪�feJ�A�ۡM2G�@��̣v"w�i]c�C!xy�����DG#����wpɱ �ƅ�4�I����_�Rl%h��<5 ������u l5�dG��&!89�U��	#W.º��)��k?i9yx2}��e𲉣�Xdt�q����B�}��p:�C�&)�F�&/[�E�Jz��..�Vと��l��I�m����	q���8O���R��ۯ^/�+�z�j�Vmm�S �Z�v�h|�;�XSqtikk��=��j>�F��%M��~ԇ�w[�2T#�h���V��B̺j1W�Z�)f��2���G�+�����ڑ�k��z5�%��;�����s(T@���!G����l&�~^�wҷ�T`RQ�"Y_�c�������P��.*&މ�}E�� �!*JJ^>>���(_��[B���㇝d���Jp�5/��Y�<��}`b�Q�����9R.�ce��8��')w��H�.6<�F���nG�xY�ۑ�g����#(�:l(���pyJ.5\��Q���}��^:��V�~��ŌMt��J�i�
-�`^_��%���]�l��ü>�[ӓ�����%��8"^7�y'�Hƭ��d����;1��:U����iN�d�O\�q�+�(>���~W��R��\��P=��+��#Ó��o�[2�?7L���j�c�?� �����bRgO��/�
�f`��m** 3Y��n:���s�x���;�XmwuFI恒�b0-��)r�W�5��W��H�7�oն�1�fA9��e(W��i���Z���8G��&D��r9)�-�඾~��Tɼ �G}@Q���-�x<=��3ʑ%���CX��o������$%���tMi:���2��i#`�N��Lё6��K��'�Р]�ﰮ��vo�Kq�=v<��6�NM\Ske|�bOͤ�U�$���8� R����+�Y.���j�4��'|`��|�^/>��o�	tQ��	I<�Y��XQb�D<[W?� ��0:�����t
b�M��2r���̒@��A�̵żS�Яƥ� ���j|�㜎Zu0�\���9gtS:+ԁ��@vUY1��]R�npmD��|'��c�+��>ix^��;a���ʖ�M{�}�,0���ы*�s%;
QO��)���Ζ`�����'`�Lע��M4�H2Ϗ\o�zv�#]q�z�[Eql:�ؙ�dq� X[!��(=�4`�PG�&�]��(�k����5}�D�f��������9krx�O�[��.N�\�k� }mj S��WE{���(��a�t/�����	�+1(�Q}�T��<1�YM��v)~��<�n���m��MɎHl�¼�l���8����`nW"�a+���J.�YEr�%Q��9��k�+h>-����[��_)��������L�z]	�niaR��$���<���t1
|O�ح���˭E�����3�#�M�W2*��@���\��z����%�Ƈ�dN�c�{��|�؉D���b�>3V��7����"(V��/Ps�`c6�恩�4��o��a�e�J��oK	�F���Z�7�%Z��X��2 'd��Zbń @�P?'r��A<�����}&��?/7@�+2�Cʓz��+آ�XY���Mzܮ��OɎ�~�Y���>W�~�:������UX��y����~@y�j���,�xP�ٵ�oK'�F�[Jz�}���x�����d%;�hJ/�8�9!i�+1�������*0������^(�Foi�U��D����31�f�6�7�ɽNM�8W�[��0K�V0{l���G�fo�Pz��A���.)! �g�3���vDfj��"!������x�tWT�ݽ�'�Hc��"���k�)|M>���0�R��d�U�bؤu�d��E����C`����vWE����UY\�ƹ�>[F���N ձ��5بݴ����UW��<���RdM<������'���߲ת*%b�Iy�PR�`�%����$i����|e���_o��蟞�'�Nx������8�A�@����"p f
||�ώf)����1+kXv�!�� �L�>��2|�B9�D���a�m3�!$�͸R�d���jSGvP��R0.=+W�11)D3�
�}�a��=%�LJ���ĹEe\�8�с�/
��L-�[x0���Y�e*��+�D�.�61�+�/㰞�>�; I�wk�^�5����ٚ�X�Z�2$�2����lZ�#(���'0��*`����D�y��k�6�
9W�wbg �� R��<#zH"u�l���U��ep%f%��Wg)QQ���B������x�����X��P4�)����ז�1e��6����Kb�|*�3!�l��I��CG"шn��c3
t5hJ��y���!�]M\���!^
���RQ�L��"�3�z�<v�f��3�,�
�Eۺ�q�7��_ٿ'�K��D�ڀ�4tF��F�9�"M���ԡ���LE�_��;���n0XʳG�y��3����GS����ݏ�4���1�a.Nv�찵;�k�g'aZNG�'9�҄SPdmKn2+��G�$�R"�ǆ�6�ӓpD`�	�~��I!6z��)J̍��qb�TUO%L|C��ef�f.��
�55H��(yWX�&3��9��{<_���ӅXsdMOkIp�C�
����|�tY�?a�m�%J1w�x�}� ��~'�#���S�����9��l7Q|���)�={�4�'�L�����R-�Z�Q�u�lDY���fC�a�2����S������K�ؠ;!u/BWI%���r�&šy�:�P��Q~��?����Bv�%���3[�L�Z�Ƽ��V��Z
���ęm�Cnx����3Z} 
M���ɕn�J�ΣА[N�
���Ʌ'�j�͠ń,׎�s���,���s;�j/ �>���	\q)�=mSXx��%�C��"�x}X��:8�G�eY��Aꨁh����dD��~һ�0q'�bE����;X���\;��Tx=�xio�2f�HďP0��nO,�����;c)%����Ć@�Ku�0J��D��8��})�Y�[��T^�	���5�~l�͋�̾>�.:!^4d��5=P ��� ���.:8��0˔����N<�^Ǳ�.��w�D Ean��ӗ`M�y���Ŗ�闡ʓ�YֿQי��m�{٢M9�<TʾNC���츩H�/8\�]�<A(�_;1@�3�5�<�AS!��Ǒ ��|L������Y���Zy�$z����O�� ���l)f����\N-�y�ݻ��(�JM�n��.���<��h�т/�H\2�/2)5��(L�!K����H1�x0���M�&���� ��!ryi4���p<��oj;��y��6��/�̮z�c�<���l�D��xﮔ����x��,jݠHI���m�f�]������Z|CgTUHK�aN���p"F1isgBH#Epq:��}��i.~�X��ۆ���D�m��
�uxDYP�^c�vbׇn����2�O��Ux�mDwO]���9�Bt�M��T4������zu%����������	?���
��Y~�����n�̦�mU��qfT� u������u�s'��2��_����s����xؼ�V&�;x0]���^��_�`:���1�G�7�FE2��>�]3�Fc�۴W�D��z�ÙZ��6ri?�*a��G�_�� j@�����gw$~���"�]�(˶=d����R:8k�IqT���V�vggg��Ài](3&d��T5em�
��R���T���y�s؁��M�)��N����I������Q
�4u���4���#U6h���Ծʭ҅Y��j/�X�2�Qֱ{��2,us6��^91K|ob��������U�U����'8�xt�Mr�J.��I�4%�#9�j�!hA6ees�����j��L*ӷ*�q`o�0�yJ��`�%Q����q��Ykj�1������dM�_םx��Z�vt.c�'�C3����X60�[S�#�A�$/�tV���̵���х5��I�oe��6�3!~W�-�O-��k��WH�trҾ<�Rʾ|�F-k~v�!�ɒ?�*�u�� �P��K�* B��#��׵9W��B�c�֖8��ӗn��[�2]AO�B���Cg��}m��R)بk�9	�A�VSd���LOD�P�h��������1[Hv��f�aDD�-�ҽY(�?3'  ���v���^}�����I�(��'��B�RD�/�O>{�~%-eV������_���w*}��b�釹(�py�����q[��H=���_\\5߅BI�,�}<��4"#�������s׶f!D���ttR�q�?I���Y��Ν;�-�|��K�R0(D�'X�֖;��!��n�$6��yb�`�?a��E5?X!��Ù���΍�-�3��e�%����Xn���(���z����D�+�������a���@���t�u��lf]�g'&tP�E&2x�=�QbX}�fhɄ$ᛸ14�^���`�-��h�����I{Z_�C.�m.�u�q?�t��3�Δ�~v���OG �S����S�G-vE�?5�9����偿҄L�̶B�1y?�3C�MY6��-���cՌLrxD�x�)�L��\^W��x�לϰ�e�f�ʊ�� ���6%x^��宯]k%��/��Q�o�ΐ/�ͫ�Ĉ�l,⧰椹݈�	q��V�s�I�fD�H��(���,ٓ��@�uI)+K��<�{@^]ⷜ�+�hr'��0B�YAh��9���sU斎�Η���'�.N�y{z�g.����1~E6+��g�5aA�4x�B�-��&�DM����4?�ޟ��x��x�e�P/�-�{�=�����+�.���ûCjS�/�ɕEg|���i&;�{�7Dt�uq#�n�Wy�?RU^q�P��<�L�w�N$1)yk�߬���spp����Vi(K��)�DXfn2P-��S?�F�����z-�ƙI�z0��ڠȚ<ƕ�J��������?z����_�keHm�LLL�g���W�������~�M�E�EK�
��3��[�[ݿ ��:��E�<��V�;��+ݻ{i��Z����������Eb�2_H&+~��dFݼgҾ̭Wx[���j���d`��o���� ����I�'�џLJ���oP�W� P	�Q�M7���>;zgZ��?L0�w�Bf O�/9)e�2��U��*�+X6o 닋ж��]�9e*Vӏ�ͱ˘��E���OlQ��>;g�4��2-δ}�_�r���5�o"]��ŭ�G���7}G_I���Y�-]7�!)��
@55p��7LFL�m�	d��II��[�����0���S�b��*Y�;[x����s��X���x�&|l���񷵵]
�6�n�h}7y��+��fhO���AZc]����y�����=8Z���P�S��T���_̑q�wm9�VcӚR�>%�[1Q�Է����7=�U͟��[�*����(�(��D��	�=�(�K����-�!V�w�w!���Q<���1����.�d-H=E#��{�0Ң�M�(ɨ�Er8!�����J�zZY�ܷ�*�~h���� �y��*h��ts�!D�VԱ-/߾��|��t�O��ݳĖ��
�Gئ&1᷶�zή��$bKj��XG��c$O��9݉Z2����\�VVݑ����M5��"��c�p,�B7έ8T�\	}�\}0��q��g$ʥזy������d�)�N ����@	bܣ��`BZ����Q�3ꅁ�M{K	6��(D����y^���2'R��6�p�k��F ~h��%�:%1��/4���3���f�cfηz�r�}HM݄N�_\8|*��K��"=,�����5X�?#� �}3T�p�_4!��<��*���t��>l{�q-�c�{\җ\������4�9H'5�ҫeV�T���h��wk��Z����0Xؠ|6�@T{5I���^�^l��v�6nx�s1.>�gd��.�i,��DI!���l:��bBB��)�MڃcdMoư�F4�(<���_��e�%����SR!�9TR�hq��D<N����c���62|�� �x������TB���IV�#_��ߛ���M�toF0�\ޢ�C�Cr2#&v���2�i�x�o$S,�蹺FN��Z�&c}�?��i���g�2�\W?>]t�Zg�i��3r���x�ˋ���|�����|G�����W�݈J�5��	��Q��}�3�	`�jo>nۍ��P���F����ռW�Ϗ3�t�xZ�¼� 洸7\�(�۷���	��w�U.���4$̥���]�%�@��̚r�\�gz'�a,��8wB���+��/K�Q���Z>�P(������O[d���N0��OP�Si�li��wtG��y���܎S��ǒ��l�Ks�:��Q�Wd?�8�0��s����TtI�+(t���#�7ؗ�I����\L�*DO�����S��,=�N7~+EG��qg���b��2}��39[�eLXzhQ��|H��乸/0I�j��3��4b���L�qF�R�x8ĹAJ�dImÓ>/�&�QK�F��jI���(�B�/�	o�(t���3�P���O:
�-JF�w�2�6*Jz�l��r[I����-:a� �cN�_�7����HCvd��꬀�Z�y�,�"�Ad|V��}����c���D���oI�+����!duoz�z"SM�gr��&�i�6�G��{AB?�ð>ksD�1�9E���;LV�a�.{2��T�.'�|q���~+�Z=N..3kk�Nӻrrr/�g��Ԁ��A�`Zt�S�R��������e��^V�h���b�#��|_�/�N��?x_��o��&^����f<^��L|g�1����&�@̞����t��4�1REǘ�DM���]K5�y��*��4Jн�]ylHǰvk"�=�Kt��]��]?Mx�\��P���N��ࡄ������N��~��7%%i��2���9[VH���J�]��HK�ʹ�ԟ��Q�ˆ�Z����|�.5�����Res~j�$�x�%ؘ=��͵������<<�_�W�$`�U'|��C�0k,�H9Nq{�PG�k��6=��<�:����5b8�N���1~S�f0��LNFi���}�ק�� /�-����½���jy�Ʉ��ʤ�͋x��D��!F�*U���$�:�h��oSih%��|rr26�3s�1�>(���t�0�g�t��g8K��D���?~{ϛ8�qx�����i=�����y$��[x{ {{6�8���un�~��}����7�X.'s�	��}q1��_�.C��=1M�Ľ������x�΋f�vG�:[l��ݤ�F��)�=���<�����G�7�/���k�v�Uq�U?�:����W����^����5i�^}�D��%0��,����K�5ھS9B Du�m�`,��?ec�ޙ?Wʠ!���E�<K�5��l?����>K�!u�K���VW�O׆�}��v�L�^���u:���ɼG�d(�%�o�u�=ǒr	�KW���,@�raƹq+i$�/;��`J��N�%�
�[�����oc,���}:���g��B3��wf+���L"0
xݘG,����ב��+fZ��� l�%Z��9���Z<V)��P����)b2�涠��nc�Is�
+g��'�o� 2�������r2�����aee%\}�A�i��EmxV���u-Q`���Q*���U����IM��K�.���|�B�d<��Ԃ�(p^h�	쐇�ƫo|Zg\����X�0�o����ӾI�$"����zq�$u��v��#|(���;�X
eLV3��_�<2��6O�9�4]��Z�L����n���;��xeܐHu��xa�X,@ս�K��휲/��{7�ǒh�*��ڦ;虚gb�Ix���o�q..�uHB�rO��R�L#��Q��]���rU��*[��ek��8�##}6��9�Ԕ�ش��VP��_��_�[0Rx����CY�a#�A�&S���U��D�U�i�P{��g�n����M�^�Y�����<�w�i���x~t#u�?�CN���d�����Z���Oj���*��+�Љ���
���1��{=��ּ��9��VyS;�=)�lB��GUC5_���������ʼfV��gE� ��\n�K;��"���L`��)�=d[����9�ܭY
,�exu���<�{�n^�\��<&���*�$�h�������?�3�zw^�8��I)1taXB��t/���T,�j
W��B�N�L�ޘeq�ȁ�alK�������/�v�>/Ϋ��B���f>3�&��^�,$?�`����x��2������v�#���,O��"l�J74nݫ<ih#x�1�������z��w˲���E��Qς��^��/��2�m1~��̊F���È]g?���ۯܒ9H�{G�#�J��|��F���Q��-S+T,Z�2)�2.�WO0����r\؈'�� ����2��g���;��x�^%:$���m\�!���ʖ}��9�o�u�s~deQ����F.�����ڐ������Ͻ<�)ꙿ?Vܜή�$O�$� '&+湓A��D5n��V7�y6��.� 6�skf�cv������R�˿+���j޾�^y�df��B�}�7qV_l�R��D<�s�S�X��JPĮl;��qՂ[��Si�=JkkU)���1@;��X罚դ����k��t`�u@tHB��J1��Q�u0���@	��(�:�7n�K��^-{�ɹx|qִ)��	؏&�1Go!��#���T���5��;�^T�W���L"ӝ��!��dxǙB��@5%EC&���O���IbԸ��|1�G�=`;���+�D�隣T�p�s���Գ�I�����;���[#-�:C|�M-=ޡj<1�yy�
�Ȗ�1bw.𥪡n����n��P��<��������b�t��9��5e����"���/�ˀ�Ve:�D(�<�{��K�J���p[�O��u1�p|�K���J��떈�e��֏���'��q���������v��t�wGI��4O�`'](�:k�q��й��9;6:������#������5�:�d��6d�X��ß �$78Q���m�k���e�����s��X��G��	�2�VT]�����9�*���z��ɒ�>�~sm��X�=��q]�3kQ����%���t��e�o�K�G���FWaX���MԜ[��
�2��8&?_�~{!JOa �����ត�go���g�FĮM�~��Ѻ�����lɛ/�8��Z�n��Kb��ީ��`���`a1��ᩚ�kJ�n��G1� ,�]#l���Հ5�f�D����"�~�[G��&����G��Y����n˗^�[�!��77"*�I���!%���l�%'t?���b��d�FEw&0��.�\{�e0�E�"\�9!'���"��KD���^����_��?��4wooAn�D��xf{D�����ͿJ�w�	�L�"���MR�0���N�9�/d��u��Q�m��DLa������;Df/}��G&� b9� _C�?��F#�q;�=���#�:=V�K���c_����1�������%�nr�+uo-�z��đ%I&����1�B��yoX�X�n�>�� 1�UB������c�'T���7�o�0]n)�W��W�nZVȗ|0���4o���r�oz6vD��H�����&O�������ԭX�2tT�k҂�;:�x�6q�l��8�䂘�;}�%Hgև0A��ջ������L���[�zDIL���[��bS3k\�M���F��4����x�)0�C�l�Zч����8!�Q"�醠	�@��뿩��r�i�A����"2��'���E�/��p�qݸ���݈���� ���#�o{ta�����Y!���v�C�f�_�<p���)򬘓e_��ޅh������5z̰�� �:?�g _�hh�����B��X�=��>���6r_'�HǓ���u-�J�=YT�C��7ɣ����n���ݜ������ׯϊ����e�]!�=�5͎W5�K2"��/�%��9^u���;�~+B`���#`Pj���r)<��\�����"�3+��J����.�P�sm�"�珹�����k4��{���qr�p�:ȱ��<��oG�P($4�:��]��:c���H����>�r(��H�7�̔����;��s 	[)d���<���Ĵk�[ގQ�|��$���pk�1��W+o���k�{�nё{_�{Z��?}-93�zu�B����ER�ʲ����3���kQ9���0�oN�����������x�Ƙ�-r������۵vPy�i.�B���w���2���5�g}k�� v�%6WSS1�( k�(v�|3rs�4�5�������^㠿��{�^�����vǢ��A�ǟ�;�y��f΢H֠� ���#�F&�=�[��l��}e˯c����\��FN��O�[�����M�v8j	����K	O&�l�| ��3+���H�������ż�/�&��p�x�4���L�}nn���}�Sf���Z< ��܆E�!� �!!!�����r��|�oa���V�є�}�u���q(�
��Sf~-�N�p,g��0���ew�#��=�$ީ4���/���J�@h����Ѩ�����$,[{VK>���=M��MR11�h�3����oI�H]>��4��&�җ�PB:�T�E=L=3��}��ЇkFW��=n�a��	���~Y�U�gV
��p<*�L7����.��4�@�=�����%4m�^���]�/��j�@��ok<u�+����FN�.�WBp��QF������gij����d�J|	��W'�����^]E�%,!��m�kr�ezV*���덑O�H8�|�J�Nվ	����;###j'���n�(�8ÕX6����%����n�3@��ތ��U�Ă�z�_�ѷ���I��u*����t&֮�Hn���Y&j��?�z��Fn�%pK,}����)�*�	��O^��q�-f��y��!2��]�\�@� �X_�';��.ĳt�'G����kg�QoHޱ��jr���S,0�40��)�᜝*��#�p<���:��Df.^����\�o�%�3ry���宧i��1�B�M�|Zv�h����ENn�\Cn�y"a�Z®^�C�;1y�Us��u��P��Ml8��l�+2�+���\*͸�I�7�́Y;�P�����PW5?��j��":�aI��hoUI�%��	��烜�����fݺ�u�"4>�=T�R���~��;W�S����\���T�ً��j*�o#����]I��Z�峪��/B"��}���"�A�V@�K7��a|�0n��8�:�Hrb�R�+��>�0�X'�֜�Ϧ�ż�<��-��V�<2��SNQ��9B]����ӞZl"Lv��rˍ��7�	�s'�v0��%44��M�tq����۷ؿ��w<��,9�X����<6.:c_��	��w�ۆ[�K�޾�'�}u�H�v����֋�������I���*�<oL�(�nѪ^�߸���Ak�R"�EI����F�Qx8.-%+::>�L�YG=���d��6~�-#���~���7#kv?(ڙ�p�B��"��d�Ԙu/mp*����n���.^�whG�����S��GSx���s�����G�#[3�
����X���w��+Tx����+�G���Ş�[�����Գ+���$T	[��=?ښ��<#���#�8�]t$�.��a�գ��(��sK[YYy��a�B�px�cll�]r�^���``��N���[�6�Q*�g��P?`��*4��6 &_��z�P��'gZ�{*�;Hld��z�彇���n;ɕ�͙FD���O���-U�Z����P�ڴ�JV�8a88�s��i3�^��hȧ�A�<V+)-a�j��2@V;-�/^���#�2��3����C�rC�[>KY�H�jsq>�8�m�i� \����ɚ/^X<R��|+��}���c����P�/>��$�P<>��k����'S�SQ&"#��������G7/�����˽)��`d+m�Qn��5O~~�=1/��sssN�����F�.��(�`�?�jI���QQ}s�IN������+��B�6�Uk�*('�Ɵ�+�H�!�������q	;G]3�����ޥ#_�f�۫���m�#n�̈Љ���a��6��:F.��׷�[�V3ic��C98JW\��Ց���Ę���@��||0��d���w�*'~u��=x𠨼8��>�<C�ޡ���IJ�����Kf7�o���^�4^	oe�q�����$٣K�K�CC�No�&*��	O�K�%���$��۽���ldD���wD>|(1��C��tތ�إ��J���&6���ZX`��Ĝ>�.�,-�����="��yf�w�
Z��㽣.�0�t���>O��=���>tq��Ue�5��n��,HQQ��#�	�T���'��t��v~_�7JHH��B��VZ#�H����#�;/f���s�"{CP�_��,���^}�͘��q�?�-��n��~:�Ǎ��}i����{�&y���ק/��d���f��~|���m�sy�-	!��.���;��r\%P;7=q_��y��/
�Ca�^�S���kI��&Q��L������C\֝��s7��N:�&ߌ����.�G��Ĺs����[�������t-�x�M�"���Ցi`u���7�HII9%~���굽n,L�ܴ���;� ���yH������S�jռGCNxj�j��+����)����Eee�����GsV�;�����������s7�<��zs�ULҧ��͇a�jjD��]������_��r� ��42rB���?�9'/�UG�^�ʍ�t�+���	r. ��.<�A�D=Wh+o��?\(��Z�H��Ŭs�
��������^w���uҁ��'E�Ȁp'//! 	$����e�pj�����������b�b:�+'��Fx�ԁ�Vp@M����_ˢ��?��K8}ݡ�~-I��߿�7qr��ǁv%�r�w8�i*7��>PMM͈;J��5�}�[㿕W>$��	�O1�f�T��aG����ÛH`��%��2�����py*���j�l��*of�W��,muu*C�aCQ���Mu����xLKۇ��N�[}�D;�+*bS�}�i��Z,FH]�������q�*@J剚���?�5��T0�I5�M���^���O�ޭ�v��=+n�`��c�z��b�g}��>i���#~���[�&M2����]7_/�{_�l��z8�ω��ɗ�4�ץ�zQ�^�Nvf�W�׌��k�p�N�*��-)�����+A��xr�	{���w}�%��.^�F����[������ ���x���^�A;��W�GԻVD=�KK�s���o+qb�׳��N��'�g���;C��'2�wi��u��3ڻO����*��U��VN��,��������#��+ģ��������]J�T���Z�2w��D����ǥ�|�OG����"Wo�p}Z��?�)q8�=���D�χ��������f���Y��Pm��R���HC�xгT^Pz�F�M�(deaD��oF�3Vb�O�^-ϧ^�嶵{���h�����I��t��y��������K�\x�ׯ��iR�{r�g�d���Q�(��7C33����������<]uXU[ӧA�)%�A$��tw��tw����t+)�]"  ���������>�W��kϚ�Ŭ9lNۅ7 2�a�u#*��:��z��0��'�\�/^0	��hY�;��5�pO��#5ൺ<ٞ�`�ۗ��ln��I�ic_�9���,��a`9؄��׋�<��!���H�H�v A�##��e��M���X:����e�[��{�`^��Ȉw==R�,:*����L0�^i�W��b�_�oAUU���}�}��Ľ0�lF�(X])�+G��@�;�քu�=���zv�"�us2i��mAw2�$��l��BGPS�7y���|P�yC��[�ؘ����֏�z.(��u�$t1㾛��֬�	p%\���ttl�/(v��e��3v�����+~=����k/o)�x�)A�G����@�ɯ:N�ƉN�ы�]]�@5m�޿��]��ݜ������M��,���,�i�=����3��Қ��O�j�0=3S3���;��fb��~y��jM#=�_�00��)�����'+��ܹ��2�������A9!Kޞ�2��&�����[UU�vrw��f)٥yi_�B�c8�� ���"��ĵ���|`�b��W5Cr
LFt*V���^�<S�:oG�<t�F�ƣ�J�@qF���N�oP����5r}XWǯ�2�Y��l���Ň��]��?�q���k"�~��32�B�j�T���+=LR�0��oɜ>����������f��U����j�QHt�(1����ܲ��>0:��F!i޷7����qF;S^���m5��}`�KM�y����d��%���`]q��#�Z�2�J��e(��<[����9��߿���C�?b�x88. �I��V_c���\�;����d���o�o�rY�nf��c޺�L}��u�O�=�툤�p����2����� 2�ꏗ����q����E�������D����_��.��t���u���-\�1���
�L��,Ȃ�@�Q��é\��,Z�f�O�����lַ�sk�����������QS�ǚ���LLKիɥ)�^]1��/�֣�k���˨=�r�M}U�K&��o~T��̛�zG��:����O&�^�_B_� �I]��<8<�q6��#R/���\!O,�crd7��Fۛ��I~����,9
)ܥ��Å �	�>VN�(���Qsފ���A
��8�ؿ��0��n��y��4a��ͩ��xNƌ&I�����닋�u��ۂI�7�s���2;z�`0����гt���?=��ҽ�}�H���m��P��ɻr׀�\��,�Җ�~��f^)S{? ��޳ǟd���{"9�������֭�6r���ˈ��#��@��Ēf4�ky!#F��^�W������(���,f����{E��+��ǂ�WuF<�Y�>	c����C���m]�d�zt�뺌?eU�Qѽ0X;����l_����I�S�W蒤Ԥ�찈���G�i�+^�냥�)�^��œ�q ���_�~B���=��5�؂<_��,(]VnK�����o�*�յ~Ʃ�we��4`����@�N�_�O1�@v��������W�Qn�/�T&v��ϫ��L6�^�B��~* 0=� ��F��HC�[J{'w̼���������P�m���R�(ϐ����<2�*8�����BN[;1C�]�q�6	��?�љڗWV6�x����s�f�Ad����|a��"����[}O�����ݚ�D1
��ee/�؁����C���ּ�<���^�5�-�JJ�I��jj���&�� ��ݎͺlk�w3+*����s�osf7s���ǉ�����`�n�'Iw쪙(�,wढ�������t}�{_�o⿑p�lmm����H{X���dX�m���&��_Y{_�$pY�$�ki���~[�헒��gdD7��pʁtQ�8��J��2zm�d�ɧܴr�Ҫ��	�hhh�>��������0k��Z�I��$>�_�[I^�L�Д���O�^��܂F*A�j&k��o'("2����5\�&J����a�K��u�dOv�Q߁J�x�L�y��r�#n��D	 �U+��O��=���s33F��2Ҙ��,���E|>��t3��5�g4�E��,��6�n��ɸ%fhH���� ^��h��F.pB�3b��Q ��D��c������^%�eI8�����p��R}��SmҚ[�`�X|R5mE�y��e�~��_n~�W}*�>�����}1�2\�=�٩Z� M���¦�p��}�Hq[��GqF����{���N+=�-��X�x�Y��2_]�g�Q`��~DӞm[{�3��,|�cJa���:V�ˋ��f��hVkn7�Jf�P�[�,�W�,s_֔��@�^�������[4��	}�K�u^�/ �1QQ���&�0�$�v�q:���_zs���-w\]]=N��'I3�N�cA���R��E4@�j�6C[�F}�y�V�����q��C���N��ީ�k����Gp�Okky��6�~���cz p.��ƅ��<�W���V�/O�g="��W;6������0�nMV������d��y�'}4_L����8,O�z�ٯ�k�v�p��|.��i{�6��$�"f��|FU���rs����<�?X�=K��1��\�@1S�C6�?��@��0����cM���������6�ܒ>�Ǐ� ����D�6bH�US��C
kj���NP�J��j]�*^�m_�=�[\���HX������jZ9m� �l�g�� ?��?o!sk���������tֻў��hd =������I�	��ht6K�b\�D�H�!4�D����X:��bz��uX�Ţɡo>O8��ܕ�������V@Pn��&��55��&�ׂ5��:(�����J�"��M�L�8C�̼<�����l!lzE��\��`N��*�`��4]�Pׅ?S�*-�7FϫZ���O<�9S��������r�c���a������ ���
�rc����i۳^�{i��B�*�9zxZ�%$���˟u��K��w�ƶ�Y�α�X[�Li�l�u����IW����^�p���Y������o���A��>�o5����9������ݻ�F��>jj�W��_rq���9�!e0e��rv�s���A�g��	�KRW�n�02�
q���vF��@�.ԙ�* )��w�9�U�zH�����#�k���}�����v�+���҃�ee�KJ^ �P� �-C�OH@���ٕ<t
�:�����V���u�зTc�p\%9�|༪���LP �b��+	�%�^Vd����Of��ā��R�٣G��VV��g�7UOv�s��� Va=��QDV��۹�x�K瞩�Rim��w�I����=��l?TQ332�ɟ�����#K7�|�+�N%��o`;��5^��p��#'Oe� ����;�yJ �P���-)qq}�L|unyl���^G�#�;��k�L�;���nt^T�9���=U}5�{��/#vbb��j�p�`�ʖ
�3t��у���������=��l��{�?<ڱgI��r�@րt�d�/�[�&��U��}av����vd������K�ތ�ɭ���7���.K	@IZMM��ժ���*_R��/AA�ㄨ@�^M�9|̄��M��Xj�m�0�Kpp��0�/�������|觔b|0�z`{hd��v�m�)v����$p)��,;0P�̂ b�<��i�G�;�Ui���-㐕���f�����hx�M���!�������T�3`�� D[�P�����zF�ӳ~0�ˑ;;��$�M�������¨~�7��Dk�EGG�T?�@�]P������� R�a``��W�	//��[i�u����	�����)99�F|s������H||ǿO[ؘ
����Fgu�k>�v�v�n����z/�WU��D}CM�=&��yW7k��z�?b����G	��z��zL�բ^靬 �*6X__���Z����;{.��I�a�-���>f�)7��:�0>&VV���U�'�߈90um8���_<���Bx�h{��k߅? îv:=+K�����*&�vyt����Z'��| �)%A<2���T9�d�$F�{��f�|�*w-...�|̮���̆N�'GA���!��3��u(㼚�zO�գԱ�읉	@�<$�v���;j��v�i��KP��<qt����T���%"�_|nAM�����4���i�cc�d@�����u��'�����WdC�)�c� ���	Xb� Y��lC�Z�ǁ���X5�d����j�J�hʂ$5+k����d��~`c`I�Cm�?Vx�^�֌o�:�]�<���U���v%앓j���Y���$,I_jQ�i�2�nMתD��D���jj��S:������M����z�.	�L�L��&͏ 3G��oQ���n��7'��4c���\\���~X�y-rw\@=x�^ }�<+˭-������aͤ]vvv&�"**��@8�R��UWZDD$+�?�+.���Z��LL
\�i؝� g^�74̀쩩�����-�Y���'mg �s,�1�j��qd�HFϞ߬$X� e�уA����wAnė;ZytD�����!k�z�'vd�����Imy�t{Fp�5�č��7���4 m'��
p��;���$K��.H��]#ʴ���)��cϹ[��1k; �v騩����n|���T�"̥44���6�R�O��%"`RקϬ�Rύ�o�hW<��4���_��<���	v�F�m��xI���uvu<�Y�5取u.�"[�w���F�����QM �f-<�K�~oPL I�_����ΪQ����đ���XЃG)K��g��=�G�W1LV��Z��[�{Dk}FB��������z!$�^m��jO���^ɻ��@��`����cٍ��t06���l� xFx�����
>&.��o�0�B�*�� �{e)�'�q����O��|-��b�yc"P�s�S��K�g�H�zA�>ٕ�����&&���z�;@��o@�4�[����|#�P�(�nY�j22�>-��j0�f�v�b$�Z::X���?�����z��C�J��vt���9�C���]�M�17R��vH�eҿ���<����Y q��2�<@���Gӹ�gĸ�m�w!�ǘ?����i�s�������BxWbW0�.}�Ch�|�US�����Cmj��1I����C���bX�'+,+p�IA�p&8��ϫul;�nm��T7)af,�&���������gʥ�l����^P����Ԣ��t�iv��}or��}� ǂP�~||���N`�����Y�l���0d$��89�������9_�ӭ�p��@�I�nLQ$7P�����.O����P�љ�P{�uV.���+�`-�hj�:=3��L]&��a��;�#y�r��Qs��J<{��Nq�9*�m-tB&j��Z��}z�?�)�;�����s�$yӛ���c��WT�\z��)Yҍ+�6x�q�Gg��B񬭿��3��8�w��
��(x��,����ܨ8��W�0ix���wm���`>�͢ckaҪȻ~d����#3��THr<��k�ۓh
(3�M�̮p#g/H8L����
�ߚ{凢1��s�Fb]d5��N\a8�.��M�_��;����cm
bd���I�S�s$�p�A�8�C]���"�i+n�AD����!�$�����mg�V����.6��}�*mT�I��w����|[MK��F�b١Vy YbX�]/QNQC�(<q��z&�XnkrB��/�����V)����}@���iϙ���m������_� a%����4th*w�]9k7iYY.T����O�� ]--) ��+�-�����X�B�����yR��z	�9$bbbm�ہL.��-�)���@��{�^�Nv�|6�Ʀ����zno��l[��H���h��hS%><2)�O� A'`z�ȸY���Ǐ�ި���R'c!�������i�cB�����?�Y��u}��}s�� ���/��9�T���0�Fׄ%%%,wg7-@�P9W`8,s/�0�.-/���'�����\�z�9۸�E��� ����9������Z/��b=�q��?3	�7)��?��22�>����u���	�i�I	0�d�G��t�z�JDћ�n�iR��۴,r�͍��\�����
�"2�׬�����C������<��U�{oL�[P��2n�r*�/"�ᛶp1���_BC�=�[L-,��Թ�0�·�f(f�!xxxf��ݾ���AD\� 9t���I����U6\���)'�n����ԔvA�B�l#��j�sE��l<�zWS����f"�LD�Bm�׊<�����{U󬸬���u�t*H�:����U�d��.[߷�OZ�Jgn=�<88��,��x����cTV�'W_�컚���4%ܴ��$a��{�~ҍ�:Z�j��W���p��r���oBQZA0\R���^p�}��*��asE>+��$\�6�"���uu�4c7.n��*""��+�և�7@�2�͜��wtw��_����V�:��!��xm�2�Ev�<`W��� ~��~���{T�(D�N��W��MD]C/���ws��&��M4@XRZ� �؁;
�$QN��5�3�6��Ѻ�<fE��](�x�ׂ�Q��x��EEC�v�a�n
j�{�'ݭ�0 ��:��͔&{`N���
��h|����'��*�N���o�\��~1��@d�
b� �r<P+"^^ۼ�{A��	��P[ʥ��گ�Jϟ��(e�p=Xr򋈌������]]��b1h!�6J[o�ܩ��~�
�������<�CJq/M���h�%�z�1[x�9a%<jt�5t3@Z$#�޷Mr!|yUU���+
zzּ���FQ�f_!�w߈�
Ld&���-��VP�ʩ�S�V��'�]Qj��Va]ˆk}i3b��z�����&���3~�G�b��*�������Ʈ�G�hH�z��0��$ɤ����\E�綞��D2b%��P�}�O�}e�uZ;;����b0S��ǊŚ���O�R����?*֔6#\9U�Ȱ/����@���--�d$��ԛ.�7������=8d"-'+�ǲ9�Q�=�*jw�mVm�QF�┨}���J�p��FԟV�.�~��(0�Iw<�?�v�'/���֏�i[Z�ψ�z8f�р���O(��x��?�k]��^u��B��ǩ�E�o�3�z�.%����������7��� .WED�ԇ�Ӎ���A�̘[��ʩ�J�Q[�� �jwkHZ�&�Ճ�u�`!E�u�쮵������%�rLB�����}�M�޴󴌲���\[�|�U}Ml)�O=���ЫPMz�Ӛ��y��R�Ƥ�Ɍץe�m;�7�]P>o���[G��|��5e��^����`F��4��3sH:��tp7��tvJ��{b��l���e�$<gd,�7}�A�뜆J,�o���)]"�젋��w�؍w#�'�1�z���((�E`��M��.�C�'�ް�fbd�ym�������t�����������۷�xx`�I�f��>����.�FiC�˼����e�� ����S�z���`�%H�v����k$=rN�K'��wK>�}� �YMf~�/�o<<S2�Z�����J�J���g֪P�o��&�쀎H:n��+�3
��i�U�l���ߣ���C��bo��q�uZ�����Ǐ������m�$�2�@�+N���B�ۋ�F�^551QQ䜜�
�\4eu�lb W�1Z�<�ĩ� +��b��l�v��J�8E���Q��^�tttL���a�JIQ	L����f��n)��}/�� �����r�� m~���8��:# n�m4܈��c�>�U�Gދy�=e���6{>�����E�9��ڮ�Q�j-@g@���{CKA�y�;�r��>��ח"�V�q�|�a;g�1Bs� ��1��,lt�d��7Q,W���yyKW���{��^W;΍T��ᖗ�-�������L���h�3��[��z�r*���uVbXD�����k��?&��f_Ub")t�6�
�v/W�s$���X�oM���� ީ9d����~D-C�u�RZw:��x������D�B��|5ž�sT=��l!�u��ݢM&��z�(M$`��,��kO���&��`����(�(+�pF�]�gb|x䄄b�5���� 4�h ��-�J�
CSqכz̽h}w-Ul[[�?������� 'k�L��TZкy|Qkgk+�W.�V���I�6Z,���>���/1�V�W~�
���6!bٜ/�L��6�w<DG���3���f�whXXzf�m���5����?�L9'1j1�B���/�Ԙ��~��DY�b�Q���D�LS@p"VV������9���9k�Q�Tv��/�$��rǨ�;���6.�1���&�L�Gkֆ�-�?�R�������s��D�i�_ܚ����m���C�H.��ga���v����r����5�Y�4����$���y����:��������o�����y��/�$Mfo&2�PͿ2�Q�9F�4K����q��9��Ñ	�c�ɟSP�rgzW�c��_�l/0*�/�SQ�N���Έ�{U�4]dj<�����)������o�Bo*B=#ѕ�>_<���(����ږPqi������'��4^ �!�Dq����2
�GZ�/4��z|��O�����.�\���]k=#�^�Nh����:������J��W�N�ù���i�?b	Uu0_�����=N�1�P�_U,`;���c3M/���F�A~�[D���C6,����
٫g�F)��]c2P��Y 񛬓95�����(ЩejG��iyT��FR!�n�ҚB��J�Mʹ�=�*�`���PRI
�`�݈��t̙�m������݄��� V�#/�t�>���W	)�M32��~;�`���>\FF��T��S�� ]�9����7����"�L畟ۭ���,TF 555�~������J�Zq{(E�j�w4��H?����2j�����q?i���.�Gv�,m�N[RΙ;:w��,@- �tt䠅vuRٸ܌JQ����&s���v�a�����E���+��t�k���1
��(��?tx�u�M��ȥ߰��MlIN��g��^F�O�����@H�}�_�RL>�q�A�.̍&�?���"u�bˆ�&kk����m��:��W1�A~����q�> K��c))�E9�\�se�@[:�kj��������j�# h��GʕSa��:��_&�5,��ߝ�}6VdP5mՅ\L4�^ϝ�)T+Խ���p�}��Qa9	M'��D=&"�w'>#�.���>W�b7;C_ұ5�����z��������X"��t�}"X�.�������������Y�����5�'Ww�gl@�W�\�~���$��M*%�����:=d��Jw�UXz:5$a_	u]|����| oh$�bascc��]0�W�>��>"��G"�ޠ�U����b�k���E��.�:w ����ٯ���%����YokFA>�������#�������ռ�k��e7��C>[Ug�Gz�ã=�o͢�d/��n��4�(���R_�4)�,��P��V�04��^�F��[>4�������}R���u�W@��O�"E1m4��m�u�Ӹ{ӄH��gَdl��/�_���=��L%� �v훚�z��`��\UWW��M&P��f!�U-�!�"؝�����N����51�Y��ۊ:�] �@��u�B�㽱/Mq�*,�I'��n�څȯ��'+,f����D���K ��6p�d�I�i�!��^�^��c�j�}�_l����&m	��c`����	p��}����+�(��@\�lQKk皮v��n�'���Ĥ��j�?j�A�Z��}�>��#�Iy�BM7��e��?�<�l~��	��wu��q"������S0х!������ݷ�_��1����-��j��H�3�`�βF����Yn�<� [���!p�% ��pt=�Ȃ���n�5��H�F�f95����^��1SV�X�{O�6�0w��IIb�y��x�����e�F�R�����f��ߕ���W����K�YXvl���g:���-��"#�7sh���m�����q��Ā͊!�͜��gt��o�C'�k�MLL�����8��v�mh#�o��յ��7=�E���I���#֎,���K�<��r�y�?~:�,x��"6*���z�E//A ��A���yyy�����u�#Z5��v���R_����6�\2�6:��k`��[���T@���帑tPV�2�o#[6eS?�g�)��;{��X7^W��m�|��T�y����aaMF�TϞ�U��Wd{�v����t��?���\X�C �ڿ`S}<��k
!�� ��Y]���l�]j�*�E�q����lz�O�>����F������H����+n�5��ci�:��v� 5WRR�d�,~F�B�͡v7�U�!�����Pf�(e�q�;�3�Y��=+�NR4�H_8���ZnN�+�a��w?�w=��߿ԩ��!� -�	y{%����A�7tp�)H
0��������#��V:1�&|�IS�Ӿ���_�x�!�����l�%��D=~1
ϗ��$yE�Z{��!�H�n����\���q���P �/�{2�1�j�e��DN�ʠȠ�� �	SaTC�q��kF���|z�Dsp��Gs��t(���r���&�ia���- ��RP��O��4$Ua5��WHh�jQ��)?���@��z2�c��$&u!֯���>t���ܬ�+���ˮ>���x��-q���P���ϱB��i���'&4���>��I�����:wx�f���l4
����1��ACEETYY9K��pUYUu���:X��i���4��C`ՃK��N,��R�k᝭2M���~����v���t��`N0�wt䄆�@�
.�|"�����9boog��7����k�� �b�UM���m���a��*Vpq�F6�X�С��ɐ���1�ݻ�#Dh��}�-�`��HT���+ ��<��CF)�M4�ϟ7YJ�<�ef���B_F*����kn]����� P��<��$X^�7�t���X��<ٻ��;�ߞpҥxD��� ����o��DGO�Pd�R^ZԹl�3�q�ۂg�z�,\ �T�sD�k�A��c �
;8�4�БJ��(����(^jzz��L����X��	L
�t,�/�ݗ��-|||������RR�w��]��ky2�wg�+N��>3����x��F#��(���/yyg�ף����Mc�a��Φ��&��#eJ�X�:��O��&U$+�����;�蓒�5�"W��A��q�3�%L7Ρw�{$��
�3:UU$�j�����G1�Nh~����;��oD�$%%��M`5^� ��;t�_����̱_ţ���
�P�J�Y��y~�a�ԯ��#��eQ勊D�)�ؔŘA�E���G�>[��_������|��S���~�b���P炞��x���N#�+����W�q��;t�� ᒞ�l��*�m�L�K4v�{�^q�l��w��0ѿ�s�NE�lG4�vP�5s+���m������R��z� ���*������ѫ7|�ZY�����,�u�}�F�Hr�f&���q��#�I�w���׮�������L�%{GPdqqq ��䕕��n��X�жs����NV/6>���&}�=o�L�g�{]�� ٚ�QPV���3:P���d�� (98<��خ/���%~��1P}�Y��c�ά0�-�G@1��Ovyg��?���Ի>PK�̼�� ��൫��C��W[9�(�<J+����s)���\�՞����N��~`�#""���bI���� 󯠠�7]�r`���}̣���R ƀP`��^�R8�sv�pB=��4� .�'S��8���0
֭F\l��m����aG��@uR��eI�Zș�1 ������m jh����/�����mП
� ș����%Y���� y��]����@(���s�R��l��h��.�F�g���-Q�G4.B�Э��ˍ�)�b��k�ww\��҅���:�l����03�������266�SyanW�M�tm�A�@>� ���>�b� �s��P�d�!l~��V�o�a� �(pg"Կ���0�uE�9��8�"8��uhh(,2R���5�wz [�'�j���Il22�.V�$�����?���!�77�]=��\���OĂM&r`@�dg�d����c�<LRԡJl�ς���Q�T�+�W�'�{zP��.���͜Cd �k쨞�t������rs��V[�������FFFP��(XP�C���^y--)##���`�,JJ��g�
Ą4�״u,��&����
hF�� T��)�ҿ�t�y��W9冞�q��%WDL�������;V���edx��]G���V&�τ�(
��w6� V�&~��y��Q���9�ql����9h��k�<>𣸂kaK��S����.r��^�|�<ldò]k0y2y��U����Eqy(�͜p;��"�!�9�
�d\\�%����o�6
��߼ѷ�2,z��*��(yC���_����9ڙN���gV��=Ą�;�����J�ؘKi}��䵬��@��&0� �|��f;��^f� $��\F����Y��x��ѝ>��4�fa	�Kq9��Σ�����#��&�bH���}�*tH��@����[��CC�DY������:s��%w�{v���,�t������~�MBWd�m�FÝ*J�'�A��C	~���uIC���w�ȦZ{�rEP�g�S��k쩖1�.��1zPn�wy���Vw��ش��fa	�5c�������ⶵ��cZJJL?�U���,/M�;� <��PK�0�O=Q"�ũs��+�f�1z�%jbB��m0��*�����A�k��|�}'`��m��ei�&�0Ar��3�
2��_`��7��,��c�jCm���Ђ�
�	�oCtX�ס���ڜ��w�!d�jj/�b�Z��(�-g2��d��F��3�>��hB	P�`�����$��N���i<��"�Y����W �)��Aj'��06�HQQQ\NNh)��n�3+55UD���Z@@�������PK��Ҳ�i�eoΛLR�w�C�n�X�?�g�;5�,�W{"�fz�A@-�����upp��(��7-�8�rtt�W��p���J��ͨ��_���q�6�����Ϫ��	]��e�e0D����\^^��ÓWU�Y��fA�$���{y�p�VS<�.W_�D�a� ��k��D��^^�����w���$X��2��ͥgbz7��	�O@��xɷo�gx�خχ�y�!x�m7��U�4�F�){OL�{FЈ�քxs���EV���I)���\*P@ K���	.���'��)�o0��bS;��kH-���]s�{�|c�����b�\�=�;C_�N�FUն����۫��ď����*�5�/�#�n���(�klr��Da��u���;6ejCh�b$!�Fޗ�lqQcg��j�����99-��^�|Y�bd����ݠW?�i���gHzz:pi�UU��yԊ��1!���Q*�hhh�4j>�kU�ũdYN�����E�U�846��4��@,�o8��Eݗ��ֻ=-��zB�O}�P�@�C�~���AܒS}�`P�U�Te�/UW>W9��]�=��dT��,��S��d��>�( �!!��ོ	o!B�)9�hHY�9�q�q=��tU2�+�\Zf>��H�U�`�ג��p�F��6��D���Ү��P6�shm0�oǇ�K7G�~�ZY��p�22�n	%&�j�}x�"�]G�#�DDz��d��.��`�m��M��6�O�}�g�1O���M/�dz^�`Wo����U�w�\�y0��������-AM���tп�}Z��F�g��IE��b�M�=C�y���4�v��[�����eb��6<���pq6�=}h S�l�d�U�Õn�<���N�(j	ū����A���j=B��f6��	1Opeڥ�����ާ.���z�LǺ̚aQQ�/■Q����)�g�T�5U�����Ufr�%"h����v}�G�I?%VВ4���>cf�-���lY�Ni�Q+��^&&&��kL>�q]�)5f 6Q�I�3u�;d7�Z�W�$]vg>e�D��5�q>Q߱��9�����.�XÉ騯�G6��4�>`'p[g�U��s=\)���z��>^�h>�8ժA��b6^B�K'�<j�r;����'*X���"~�п�ɥ��Ǯ(?��4++�	��RKW�5N�{�N�SV�$p���������I	�]}���Z):�����h�;>CS��_*��=㦶�n@�B�0$ᲀ�x��`�����͒%�q��$����P�r��9x�V�j��]���e���\�aʎz)w8�z7��DwL
�3���Q?~P
^n���p�:mO,-/+��3lI�P*�����D�Ԥ[��T���aE��OA�j�����=���=ի{ͨo�Gu�j���<���2�b��|E���4P�j�+6������}U�	�ّ#��3��'��j�/Rs_Qv�A���T��"��h����\����.7�������%��#���84C5�CZMJ��W�^��;ߜ�b�.�=���{���Ǭ�E��m��v���Nb�vT�OA'�]�E �9?$��t?�Q8?N��3Y��֙��nI'���\z8^'�����Ӕ�懾Tx�]Үp1r�� bV�@h@�T��Fu�*�U�����1�[D��$:������v����N��y,�ەӲ��F[�ni�E�zT:��eU�:���UN�_t8��/�
�(��(���r=�A�C��SH����NXM{�Q���̻�W:��s�ԙr�#���o9#�>��z�sns�3��DX�K����[�����b�Y1�(���xv���>�U�1h�.�x��S��(�#U�t>'+y!޼0-;���[(Q㠱������3t@���v(ڌ����grp��ծvooXz��;>����7�r{���Q\�.�~T(��ᗷ��|PՄNʉ��sYMhA%^�1��.�=�&E�S����Տ
j��4�g������L�K�� �h�6U��uu�&/u��5�b���Z`hͳz%S Ή����Y� �7~wE_���������xc)a�3���N
��^��|-�jP�O�W�	��Mo�\�����-���%����懩*v �r�^הR��׷�P��O�,��5;�FZBd�2���
�c[�쓂�"�L�PW��f���jU(��lOFZ��Q֔��6�:������᜴�OS{����|^̲?d�^���ؖx���'j	��c��-�1`�
�fa���t�8�sV�W�yA���d����,0PQ�1�4~�GDI��ĵa�WT
$A�hE�C^�N ��YΧi *ޅ�[CCR�˽<zrM����.��\~��T�Kx3�9O������	ܫZ֋�~���޺v��$��4ۜ�_�j\�}�|>g|���Ϝ���O�ɒM�z�) J���뼶)@%��X��>��	�,;?�����-b�0#���F:�������A�.�-��ր�����i깡��D��T�`�3��p�y�;&��T��}�>Wٔ�7>�<�
�����yH瓳7m*F����iA�H���u,76�]�ng�g�c�I�P2j�۱��h�l�W�|V-�%��̖Bo��0���Lz�ȿd3��8Rs��$��
'��g$�5�F'd�ji1�n�ɿ'lU��
�E��M�O
|!(7�g 6��h`u���������z��'u�p��r�ڂ�����x�&�Qt�%<_� �D �u��4̬vM0?�mb���OBe&�K�A�^��z�sh�W��sT�%S�j�,H�����{�\}:&��'�"�-]R_X���ub\�g���OCX�>�`���N����&D�.�D(�A��9.X5�r�������Ĵ���,|������0I�;���4|�� ���Q����?8/uMq��o��L�)��3ǎ�\�أ�!ɗ���)�O�(��s�ݕ����Tp�k�t�	�n���gG�����H��~�Rx4��-y��U`�f>�[���"X;a,���b�����B�$%����\:�QI�6�n�a�E-%�@��t���e�0wWZ�ԯhR�J�޳���7!~�N��L��6��k󔤤�=����j��16�8>G��'R/�%���T�N�4I�4V�!��j0���Y��^~{��H���5���<�}_��mؐ��6�����F���J�Ke#N��/�&��N���BXcF��0�~��`�k���Ѳ���Y��#^��o߾�L@iz}��޴��_�т�l�G�B:x�Ѓ�	���.�PcPp�^�z�j�v�[z	*�Dh�H:9��%	WH<<}��栃ξ��P��i{H*H2���K6'=X��IXR���@`���,���d�g�j��4 �a���u}2�ۮ-|[���w�Ys�R�Q���X��VW�Iz๬g�}���4���zVWuw��k�.��N��%\��(S��(�U�Ua>�8s }Ax��Ԇ˭g�K�S�[&+��OM/V�ʸa*����kd'W��4s1>�S��k��4���~�]�
���z}���x������($��Y�������l�wYWc�B����=T�u$�Wp�3������l0����vH��)�e4��RP)\�Z0ay?�����Y
������������iL�+�	����C7qS��duu�[zH���e��.��Ύ-l��R��8d��@�E�1�n�@JĨ�S0WԴA�1�3K�c�T�����g�0���q��7�D^ �,����
������fg�B�΃�;�g׀'�!^ǔ�E)w�(�j��$�Z�'Z�V̹@7C#5P>���ۂj�_G[��u��bN}Y)�d$Yl�4��qL"�*�	��%�Ѭ��U������w�m�
e��^��i�r�J�]y=��(�BW��'�i>����-��Yb�U�s��2���)����E����H��|@�/7��O�'�&p�2�شn�dx�U�q�-��[a9{���6-����d�y��%hp�k�Z���Vׁw�Z�`)�𻾻gʫ�W1�&�(S�m��[�7e����6޴.��.q���B|������Cq�'�͹� ��K�w�2"f���_���ǡ�h��w#y�
����RT"�I�����8�@��x7��9]��{I� �zl�gv��1�f��+�}t)K#�V��R�M���B��z���_{_����=cƖ%ɚ=cK��-�Ƅ���|l�}��K�	��Lv�d�l�G"dɾ�,�������y����o�׼�^�}�s������s_�>�FA���_}Ť��1U��}ً�V�	]y��9�rn�B0ܡ��"���^��&I�����ϰ�	r����<�>�"wP���f�h9Ǟ��\��� �vuBB0�1�Y�9U�k?{�ڪG���^�-�O\����=���9:�����>���^�����An�U,��5���p��w�պ���'g|E��e>I.~:����x�p9����!��7���2L��'�ᩥ���s����ഉഋf�"*�ZX��?x�B��峓]�88nN�rP�������@Y���\t;K!����ݢإ7g8����_J
�I�ٕs���~������̯��l��
�Ƈ���%}vO|���X��l�4W.6I�hO��k,���E�*�ە��QTNK�9��1E��O�юг� ��E�����I�E�3�8�ܺJsH`C�``<e{i;Z��Z�x !�3d�ƦˁI.7)�p�cض�������%p�kp�U�����\
��*�Mv�ū���/���Ґ>Z�qٛ�Z4�H"9���3E����	��V=��(�\�LM�=�.��3�����Ժ�of*F����n99޸E�S	���1} 4E�I���[k��YX�šL6=����+avNP'��˕ӗ~4����h6
���:d��vn2t����mP������}�n�;��������~0������>M���ӷj�.I7�5mx�����B�N�V^�e�2k�N.�U�ER�X�$�-����f�j��rt�o2��O�DZ��4.������m�:�.,-m��MR=9�V�\8�2Q#�j���^�+����܃k�Vڠ�I�6y]���'h���ŭ���^y������L�L>��[�bL5r�ZWd�!WB#�������P�c����	�[P���^�ͪ�=н��l���3ŭOIz佖�,F�U݁i�\܊�5+��&h��[X\�d����`��H�JP"�_ID�F �jb�31��n���}+<�ƀ�O�4"�v�

����؉08by�A���k����_N�Bq)y
��hP��P�2&��p����F�[�����_��ӂ܁�
-���5_���gu'Q��n����(@�oob���7魺�[Z���vE����\uC�X�|0R~;[>�1'8ub�C�a�э(�Yt2�A�0���_���E�4f�/H�+dH��0+X��B�/:$]���y������`�����A�P������]���L��#p=��9�b�p�wW��/��?�F�"�ѳ x�|@a���Z�����}����%�K���� �7�ti0]�:����!�����|y��@�E@��:t��m 1}m���V����e]�<��Qo�&%�j��AX��d�3�?$dff�;Ja�����K��������-G��Xe��/F�e��MǑa�HF�fq);;�/�����8�ii�6��H ]*t-�<�ɮ��ydڦ�M�Rl�px�͡W��������&�?���$[vvu�|z$쿓xKB\|��	 ��AA@�L�!� �v^`�Ri{^[�-�R�����0좬�ZޟnT�C�|�!����50F���p,����L�ņ%[D�\ziA�mc�p_�hZ��N�lQ��"���p��rn�yg=B�jY��.$���f]���S=�]"ў���J�S�3 -,yĶ/����M/�����:7� 
�*�r�-O��SE�z eĀ#�����$���5�mq��2�0����dilq�)��@	1�h�^L�-���:�<�s�$��.����^N��YIF�FT�DTm��U##��EO��<�R��~����+,բ�����c>���6��G�K���g�cB9p�s���2���t|��ݕ'@rAG�ǫ��(*j�6�͊������
n�%s8(�c07y�6t3!oz5��n�Z5)�% �Wx��gN]Ǩ�����?��i��.���,����"�!Ҟ	�ݨI"�f���22���o��x�B��J�����l+�Ұ�'��{�QB�ȕ�Zup|=8}Ӧ,��\@�AP|{E�m!�2v~N]���.�������z�8�0��4�������#���`8���tՍ�Y�	��֭q�&���zV zzA��c9P*^�>Ev�z3�Zh����|&W��2֩�H;�م���+� b����C�Cۇ~�qP���ȫ���s�ܑ��~D[]�{k����)	̵cH4d���"�������Q�A���H���h0���r<EH�����o�Z��@- �<;|���NWy�=t��pLwh�r<fK�Z㦿V\KM�u�>�i�=�vf7�'Q�r)W,����]3z�s�l(�p�E=���]b�v c���ӥ�54V�m��(X��3U`�~��!
�(i�a�3>a��9߬Δ�չ��7��H��a��/�O_z����r<�i%��<�V(R�\(2N�o�ʣ�b��wxp7@�-��RR��f����i�޿}��~���$��cPO�Y�)�����t��N�O��P�����I����yŧ*�_0����}1� !8�����@�.fK@��|/`�/���~�Х�w��M����H:�$����s_¤�.4]'�#}{l����ܫ*`��H��Up�Ӟ��t��/ϲ�c�"� U���Ϳmc�N`�OS��.���������;A0��z�d���Z!�l
؜�����=K]�6u_�11QZ���gY1�MI���8K�e���ѯ��R�tPuaa�a��h~��p(��=EA�^�vK�Гo��X�+�|@�W;�I�����G�
٩үZ��a� J�����@djvj庮�ONZ��-YDe)�){��n/0�����!�����QAwY{܅I3�c�A�*����%�I�W������::
��h�i�2ف��5�{�`�6CD��b'[v{�M6t\�8R�=$<�y]�2�z�Ҧ�+�4��{�2�؂�gysWXWu�z�� ��!�)�:�oԭl�dC��?�R�M[!���
iq�`ླྀ���s�d��~�u�*?�Օh8��Z���l����.GD%��I6��P��վT�a�A8���`�	���F�S�@����Ia��V�Y\�"W���g�m鹙�`�ڴ>+O����N2�dۯ9ӋfU��!"X�\@�3e�H�s� a���bC�{4��o�@pD���1d��b�z��SSS���ύw�m���El� �/�Z�(v����Cxw��	�ba'#B��G�2���C���9��FO�D��7�4L�՘E��A�6z.�䦆��^�l+#��j���x��]�Q�A
Z��P(�c�Т��d�T����V?E�c��p��x�b
3o�Jn��:PY3��+�L��ôM�y��ɷ�;��ב�GCN�9z�gu��M�"�	�g���^=iN�ru� ��v�Ս~4����פ�.��pwm�d�o��Gz u���2���`j�QI�g��8��6��V:dmuAT�{!&_j^+M�)�4f�������b�e�jL�ial}��vQ�}0��!�?�(�gaV��{�|^�B��wT�mIS��(Z�蠕����
=�O�#V�n���s�-4�%���r�<9��i�V{�F8��vOk�Dڗ�����wɋ�.��|�xS���h�_���U/3���_Ш��Z����E�LX��"�pND$�2��6���ԕC��E�~�菞�1�� ��C��8�4#�LH�t��V��Q<�X��zԚ�LJX	.R�ZH�w�v�v&���x�O}	څ�O�w�ec�6��5���`v6fr~~��pZ�%�U/����©s�Ր�5{����#��j��@i/�zx��H���񢏎�1G�6��|�$"��]ow|��x�kC�K}�f�
IҪ����'���5ގ J`̛Ncu��Ĩ7]'j��}�Q���N�v�rh�� ��p[4oOh��~^�P7k��@�'pMm�\	��t��f�vܑ�;�W�W�|~є�g�2.e^s�J�+�Zh�K�]��4Ew����W~؃�E<M|���F��6ºu+~"	�;/��! C�3�73��!蔹���
�]��cj�
ZO�N������|�TIc�J@<!;}�$!�� 1+��p���Q���R�JA��L.��>ƨz�$��6�D��"�k��5��O7��(��'�M�UŞ�	W���2Q�>�Y�����R	<�� �%����f �&��˅�_��VC*�ؚs]ޯ�k=U�m��)>dG�(ˠ�)_�)�Ͱݵ�E��O�MWX�����f��W����t��9C�n�X�̔�JO��'L������w'`f��n|�[�*Ny��Y��b8Ր/���[�1:`o�+(r:I�:�+B9�=�}ȟ�,F�HI�'~Zdfv��U]X ��P���2��P�qAKC2(����S7�����)v�] :@�������?\�>�8:x-FC�&1{i=)�>0[���~փ���� �0��k�R��G�Y�gto�����vJ���
�t�ƍo-�\����gN��L�(6�-e�?X�)���2��Z�Y+�1���RS�;���dY?��J�)))76���?Í�-���$+�?��M�b�%��C���w�n���A�Մ�+E�J��m��2���쫓C���J"����
�e��D�dL��!}���>�ޝ�m�-�	m!�nEsoܤ�Qt+p��o/�j�D��c��iy�:p6�Ɖ�J�I�X��o��W�H-�*��?HEy��8��y*",�Y�_�sOW���l׏��G�_�Z�1-U�@��rv�����g#W�5Ѫ��׺�?s��Alӧ�eq�Q���ڄq ��6�4�t48���=|ǋI�J^c��sF(����b�{C���T�0��2>��@��݊�<��8 �nS��H���R�T� }�x`$sf�b����%�P_�Q��%����-ܴ�<�t�(�X�-ƇE�vvv��P4��>~���J1����h�4�Jk��)Rt ����J^���Ԡ�3J1(u�Y���r��RS���=� ������Y~�sY~3s�O�CJ�ź q�nS�߫y@*�Ag�ా��ɺu�ޒ���� Nb�A�_ݰ��e�-EQ���`R���$]'!9���&��<
.�m��/6��; �o�����R3��P˝�o��j^�V��7w��ϐ1B�Dki�:ɑ�[���`���jM�r�t��.���߾W�� �_- y8���G 6�c���Ҡ���V͍�[h%��f(����󹪀j^noQB���U��.�H���C[  �"��gKR�9���2Q�g�9�ش~���
����wh%¾�ϯ�m � �67��7;��6����hK����^5�R_����ۤ�UΪ�՟��9�*�o�5���Q)��FDc���Z%�}��m B�o�tN~��u0�5�h����8B?���r��7�f�.A5zr����b��C��EO�6!1�]�^-����P�
X�I�'v `6Ж�}��6�>ӎh��2|f��N���d����͏�8Ж=b9A�b�m6��|�=����+m��A�p9>�{��  ��Zw�f>Ȍ��ZP�Tf~J��Yes�wy;�F�	��T�Ԥ�pZd-�2�v��;�q�������A�e?�l|և9��
�)�#��Yч&wk�+��B�*��B�ʃ��#�{��� P����M�㺛��k١�C��!��IIg�،t�$XTOj��#���?�!�b���ݾw�����jP�߹�ɂ������-���r��y9��_0K֏8u�o��kMS�����B7k7�=���C	�����Io�pD�jE[C1W�?{�E�j� ��߀��v4.�85��*��Y�}�h�E�0�)i���ŭ��4]%!eV%�8:o�Ҵ�N��H����Y���SyY
@��)'L�������c7nz�>��:Hn�C%�bbљ��� jmL7��g�5m
������XjQG����h��I�b��7� �9>�3�9aPE>�,`���n>�?�O����k��(�G��KWt���.���'<>,��Qr�A� �i'	Jc!M��p;%�	Y�����ʗ�)Ö��pL�}���O�u|-�:��6U����dd�h7�R�ʨ���qp�9�^a�g37b�	~v��k�z{������G��.��mQL�����d����Jc=ah�O	����<�,DT�*ɺ4�߉sN-�G�4��5���*3�����7Pp����xvٽ�XZa^���6�b30x��ƍPǫ����g<_>��W=��f��}��]3+����Ӫk[YY��"���3��2sb\��p!(v���J��V�Pspx���F���X* n���S�ډ�<zs3t����h����'�<��GȆ� _������[�ƴ<Ƚ��������$��tC>I�%u�ֹzbpɠqp�ZD(g�w����]�}U�e�k��3P���o��m�uI"q�E�8$�N&�Ӧ��g�uS��0�ȴ��PW,C|�<w����U7�m��eIq�I�� t`՜9j���]�Z���V�X.��yG�i�@���@��!!��L��CΈgafl��>�C�B�w��5�#bħ�]iǵ��x��L�(*�W�'Ǚ�[�u��1�~���
�h�����r�]eL����>�BȪc6�G�Ŵ�6����j���K� -}�@�t�3ԝk��QJ@a	(��i��-�%��^����?$p8���/��}�d������ ����o���AR�	w�Jj�|��H��|�Z�(����FQ��qY��W���q��x\=-�R�؆�{���n`��@���q��/���*Ը�p[�xk�m�����`���%p}���bL=z�����u[cB���7�	P+�]���[�Wn԰�IL}8~�h���S���cp����=���l��[ׄ��]��d�	�R�UL�����Y����K�7N��oJ/A�p�߼Y��&P��6�U� �2�|�.d�u���u���ۏ8�/�b�K�zz�P���>�������ҷ�]��<�t���bt�����l;>��+J���c1c:R^�h�~��h�������0�[S��g�o���<���ƥ���~���l���Y��TQT=�I$e.O�P��.}āp��ա"���ɴ�,ȥ��!�`��=|�l�i���ߠ -�SPY�!�40��2���{�҃�LS��4�jg<cϳ���L�1��L4؏�ǐ�̬���?���c���O7)��ur!G�����p��SVuX�����lt1�r��$]�w���M�R��_��H�<��(t^R���o�]�{+�NV�`��@����.t�|�m�L�#����2�%f��J�qr����)�WQ�m��Ȃ�e3v��52�M˄,������)��
��\WX����[���6J�t���U�HA.pՎ�de�+���i��<U�&�pf�HtFfil���3Q�;�%�)Oa֫el�k*���|��iĬ�[���DM�L�����1��e����������װ�6��ƬCz�(�-D���$�&���G��u(���RNhH��0j��Ʈ������E�6Z1��������*�z�dhst��O�o�1���ueA��*i�9�H*��zpM��24���=:�9Y��BՋ�>M�ض�M��h�oȦY���|���m��nX��+���z�e3q����{���u��PK   ��{XF&�!    /   images/24a54a69-5cbe-4d66-9ad9-6bf107554def.png��PNG

   IHDR   d   (   x_C   	pHYs  b�  b�<2�   tEXtSoftware www.inkscape.org��<  �IDATx��[	t\Wy�޼�wI3�,Y�%y����=!N�Ҕ�@Yþ�@��ۡ,'
(phiI�B
	�,l	Y��N�cǋ$[�dY�H�h���w�{��Hr�=�=\{4o޼w߽��}��c��kU44M���'�j�ڝUT+���������^�Tas���ɇ�]C,_����R	6���Kv��h��׼��x�"���Bk0,Ǖ�@5�Mtd�WD���(s���|<�`S��6�����*ʕUzWͩ�d�T��o�8�r	�NM"/£�f������9�e܍��舆�v�".y�L
sM����<�6�D6��n��8�U
��{�.�|>T��5ݎR����
���f�[�Ē��bĢ�r:�TH!d���9"�7�V�A��¶�!�z�P8���ũX�փ��f�r�g�bGE!m!7ڃ��
�v;�J �q`C��3S(����� B��~|'q�=w�vJ��"����c|���lN����}���e!�����H�.HaC�'&sx��V�=�������J�jr2B�EY���,�g4�x���h��J��躆���r�)umc��Y�F�����c�M�R�M��Ahʦ�KY�h6mU�۴e+g?<���D��ʰkeL�C.�EI�hw�#^tb� O&VxQI���Ɇ>p�:_q8�y�KI���ྜྷ���Cb��?S!l6����$���߹i�z���4e!N�o������y?���֗���!�.���!�/���|� ��R\T�`�!�����f���xd�l	99��+��D�\	��&�>�]��s��8u�^;S���R$E_Z����v���+eԷb��d��_ن�~�=H����Gvߌ{㽈�X��ē���N%Q�W��lw�en
�z{\^�p}��ʕ�jZ����)���~�llCFa��g��C������/��JMȗe�Rgoc�X�T8U*����)�R��a(�m��C�2��L)�R�2ƿ��w?>���K*�\�=*�?%�s�����x�E/�/�g����i5�t.��+�p�x��8q˔(v4G�b��|��c� )��(�W仂r�2΄x�C�d�!�!���2h��6���e���7ee��?����H�((.͍!37���Eo���놌�]]����y���4k$F5(Q�o��U�q�m*<�d �^����#�;hL6[<5�ΫdK���C9w�ǲh]c�A1��X�E������??���o�F���Wu�I�A��xW�+�JE<�lF<ځ��)���s�Kn��A&�2��JX1��]�ӋiL	4#��5�ʂ8|Ϊ�lˍ�U�A�t�eMi
��K��_K?�~��ى��s!L�9W��C(�k��ta9�Rr�ƾ|}J�����,�N"��ڜ���P�,�q���t+O��nE�9I��U��-���r��t�^r-���÷8_�uV���W`�D���s��%��Ĩ�~\%Z������Ԅ�E/��4�A�
�%���G�Ђ~��\��Fx���]yň���B�|���x�jZm�e�Ǎ�[�oL�얹�m��F�G%4���h&v�Ӂx���ہ�&��bY�m���J���:���߂͏�)��d�?���t�J��������pߊI�(K�W�?�7��b�$P)v�J��o�v��w�@*FΑ�U�eX��^���,e��\���<���R��xs����xow�Oy����<��RV�?йC�I��m�����M��,~|�����pud�EbI8l�`���o��aA+�P�\�����=3�}�x����������9����ۿC�+b����A3���+D�g�~�ʋ�06���̪<�6�
8L��	J+!�++%POk���F��o���x���!1�ο��q�bT��j��y�s��A|��sQ��h�y�4�G�'���u�m�M(e4�F=K,~��12q.���{a+	�v�����6^�c�V5xBO����־��'6�H)��( ޷uc�i���\X4�q��e�Td�����v�I���b��1��s(���$RL$/�ExeAe^�3t5��*���ma8�N<u���;�حrqE�[X��%7|B�]4�ʁ��r˚϶+��Π
�%�E��P�����X�[�R0��	��D�g��V	�6<3����N"�+��U��#8>�Ɓ�Zh�Xv�Ex��$�li�=O��Z���2*!{���r��&���)K���w�a��y�K7�c�� �F�W��0���v?�=���o�,�L%�Q=�m��^E�	�.,�6��񂳺�wd�d�qQ�[�mEH��t�����ozu��m���]#;� b�C��6����c52����\�o�H��3�>���56�q[�$QqY�L���܁��_�A�zZT2ط��5�P�F�ǰ����7Q`II��h��5)�8ω�)C�2���?���Η����q9�RF�幃�B4�9��W�丢cx6�8��ɸ
VTa�\�q���6��7�T�O��]�зi���"��E=౽��~
[XW!��^�έ�I�vU�2�nU����B]���^7
(p�.�j$y���9���s۱�ţ�+{Ԅ8�M~|�W�+��NJ`� ��^
����w���o����q����G�����R�G����Ŝ�� �~�"��d�6��cGwX�\�KP��LJ1�M�5/y��Sh�GW%Mq������WF��|���q�p�K^S�-,|tKSeB�k���
��Cm�h�ގT|���a�E��	_0�2!ʨt}ZsG��]؉C�I�f�y��Ds"��!�� 
��ꪳ[�2�ˤF廌$v)�OK�WY^�w�E�?�ǧ,��ŭ�pL,��݇��w��qَ(^�{�T:J&O����vpz!'B/���"�`QP�S�:��#���e�$�y_�$�(&2Fq��f|9I�;\�ގ��A���B.����������?}�ե񝑵�'�*�Й����p���R?:$I��Z����c,t��C箉�:~`��&uwCR%<|h~ER����O��M�U�g��=�W̻�k�F�hk2�07����}e�O���xB}��ߌ�B�ED:?{�&cYl����*��[��Y6y��p�CbxL�?��#7x� ��Ղ#�x��r�>�O�㫮��}$1��}��n������e]�q��!~���|x}^e�|�/J⃟��}aD:�V߬��1{\���n��z�ۈ�?S
��H��bh�G��ݶ����K���g�"g�3�]T��f�#�o4s�T�ݶiR)csi�Qh���2�nd�Ud� �q�Exۋ���s��z�>��ݡ*�,�|8�\%+Z����+�CYց*���R!?̌���mp�=�~�a��>|� ���{��ij�<���,�b������;3��L��ϖ����ZH3�56��n�>����S����`[V�zVd�s+��tw�s���gdC�~ 6�^���ۛQ�d���W���h4҃c����O�������O~�������{qe�.��z_5P(�r�%J�B��~�"��%�A6����:�o�+�Y���^�%��(�sJ(�L��*-�jb����=	/6�o� �BP��D^6����h��^ANEU4�e[Be-A'�Kn�U�\��p�'�b�a	���D����B���C��:?�Ų��<�~�@6��T��\H#�/�N����Ai8,�fr�T\Nˣ�2�hȋ���q���������5/{6���\����/������"=�}�Nv�����l��Yxͩ�a��l�e�R��Y���pɂ���x(t�Y��0�	�K�`�u�uc�MbZIA�>�Md�Is�cr>��TA�v��x�s��k�TQр�����Y�k7J"�cB:9w��5�%QsB�O�j�R>'���h��ʠ���,~��^��|a���BL)��M=H�O�u��XE��y�~�P^w�V|��'�-(���a�FSLL��zH��KHrOIL�Ġۍ|&_�Fd���o$E�|�_�f�'̜�E����;�Ea	�
�E�G!�s8�rÚ����u\b�D���]�G29%ON�6�l�<kJJ/���s
b~AVY%�&>;]D}	�^�U�2�+���+77����8KE�y���<�kU$S���/o���k�؜�뾵��=!����{�w��c�9�$��k���~7ԏP8P�ɱ�8��'в�ê�b�l@`kD-���l
�R֜(tza0?#��C$CG+��˪.L�
b#�g�8�!��@O��*�00�{�xì=��G�� �v.�S�wl*��HJf5/,�̏fːˏ�bŌ
��S�I���gjƿ��x�^Qc�������sNq�������,�[I�����lƩ���?�5��)�8���2��w���g��"Ǒ4W�&a kǆ��HƬ�c
�|��-Te�ԯBX�UR�lϞL.�A`X2���)AY|W�̌%\�	,y��(�M��B{n3���?:�E4�R�9:�X1��|ȹx��u[)<.�%�2���<� a��'Yi���r�ӉC(]��ׂ�%��ᮔRa��r�VHF�j���B�!-h�c�ZT���ju͐al�����^#Q�϶�?[�3�w&xP���1��/%�qۃv����vy���� ���`Fo��Q�m�+_�
��v8]nu��^��ϋf�rW�d�W�z_prK�)�q���B[y2�H�VT�+�ڻ��2��@�q�UW&k����#bqDE<��Ev��F���a�nai�01�D�|d���5�A�c�b.�
�V�d٤IP�B�R�=�KƐ��R}L�/?3��+�V(�6�UW��&�#b[^=�ࢋ�F��K��O_����YMVW/����3C'�>t+���-g��b�(.�~׷�X�\�;�������k!�{CxD�u�
�bU]Qc��|E��`��&���B1��`��$o�`����nlI!:
���j.�F�)�&
�5�R*js�R�<����R����Z����\��_\ʋB�I)Cao@���'�%��{6���Or�xJ)-֩���Ǧ�/.J8�v�[1t�kTaQ��Q�*��"�#��U��V�?�`l~S�=��J���0�s����p"�����y�[�(kK����b��[�BYDh�>BY�3�ד>��(��������bC>Yq|\s�Y̫�&�����ěox8�ǰ�݃��r&/�oy��[\ʩ5��d1ּ�,:����W����n\r���Ó󯻲�8�)i��g7������h��ԉ��X8�O�S�'�h��j��\⎓ʺd�VOp;4U����!�,��zU�J�'t����k�S��x���č�B�@�!�:a/C	�jSU���1d)���2#�3I��x&2|���:���m���2��o�AQ�m�i�OZ�{t�`��pv��(/�T���Z�

S����;�?�O{����v���~Qt��/�~��mh���8���%ƛ�G���k�N�c*�%'�����e�fNY.�Na�1���^PB#��gc	Զ��N럊�B��?����pʗ�!�|H*IYT��u��T.���7҅$����;V�2��&�`��|聉E�q|QW}c?�b)�K.r�;:��e���]�gdZr���� ~r��V�B(kl�d(;�(.
݇O}�RUl,ˀw�e�U�e������-]kj�ڥB��)~R������q������eȝ�wg�(����C!��l��א2%�����U�d^�K�(��w�Q���uv�*�dב��;������jwesĂ���ϕB��|<8!1?]W�#۔$4y/��IjZB�����.�sx������Zs�Us�dhm��3����
���n�R̈́���Z�ʺ�RD��,"i%��v!k����z�d|�SD]1��5R�;���Kv��KBse%t0>��WU�3)��>���N���.��DoK--���3�QY����F�`����0������C�n	�0�!����G\����91������7BW�sk֮�p�0E���\6�VEU%Aq�_�~�dB��-��Y'���eX�ξ�R
� ��"ب�6��"d$���ߞ7��\��<tr^�ۻ��@u��8.C'V���=/� ����0�O���t�woEh���{xa]�)���v�@�ԕ+fu�*�:	[S�X�Dfn�rzBpx�
S \�"�dlg��Be���*�ֻ�j#���k�կ��<'�dQy%w�̘�iA`�˪29�1�lmcj�6���H�˵}�:����!-���'T�h-$��=��rV�VC�^FUľ�%������A�L�a�C��*�!f�^q�x���it��b�̀�a�3�^�O̧���[U�Ya�tOMbt1��cs��߮���܂&��i�ы�@�|&w0
��s�"�LkeY��#1���.$:�Y��+�U�ʫ�@^E�
��p���>W[Sۛ<ʺYBo�d���I�^G�c!7֫���ښa]v�o�`���饄�E��
�^�{�{ў�DE#�p ���$�e1��W`C+�˿���	���f�:��>&Qe3���8��|�ׇ�%Z�h��z�A���J|�_��������&c��\7z�4n�um�{���Q˪*�[Q�0V2�P���K[�`�T9���~��0��
�}������2����[��E��|�"G����*��9L��0��ᩔ*8��{,q��28T}h7��J�*��֌�ebsr��4�_������^�Z�Ru
���ƻq@&5]x7���۰{gQ7�Ne��� �;��pd�'�K���8��Fx뷔@��&n����E'2g�#6G+�:<��B%������B[��ϛ;HXza���F��G��N/<8�Tװ���%��R%�bņ�g/���5c��¡��1�IG/�Z)�
ɠ�J(��zQ�*pWBH���t�v�7��L��Et���|�����\��w���T���4S����Q�Le��2a	�/J�{��um���΀�	a�d��	7m����Se������A��B3yKm�X����9�(ֲ(x&x�>��h�Z}L��|����.^��!��2p[��\�
�O�,fʹ���s1�yX>��*��%�c���4\�3�+Y��f��n)�5!��D����3W�dW�.�o�H�7�~tZmAP��TC<������2�\-T��Jyrt^��w�S��~+��-���c�;�{�de��b�;�vr]�Xߑ?{���X_ɻN��ŵtc=���Y,#��1��1����߸&2K ��&���A2pE-w)_l���C*�T��L�w�B8���S��ڌUAqkw&RYL>���ƅ��?$Z���X�y��fZ���bx<�.1��4҅��s����E~��63    IEND�B`�PK   ���X��g� 
  �	  /   images/4f5a6b59-a216-44d1-a198-112719b334c8.png�	��PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��ZkLTG�e���	>*���M����ZMl����iҪi��j[�?jb�c���X�hml��1��b�A� � >A�
"�"����;8ܽ�h�Bz�q�;��>gf��^�'OV�a�i�b�}v�?^���W*���{`�
� X/��У
���			���Ǣ��M<y�DX,���,����v�_�GL�����1bĈ���^o�~εZ����E�l6QQQ!z��B/^,���E^^�=&&&J���������GDD�N�0��# ��[�n�:�N{0E]A|		�� ������q�ƉK�.��[\\�p8�Ff=�x��SSS#��;��YWW��1YYY<x��������@pa�$�LNNv��+�j��@��ӧO[\\�i����;`Ȑ!b���F%y4�KyR�w����o�����;�P����ݻ-Z�r��=QYY)`���ŋ�B<�����3��*CQ7>kt���h�th	�������?��ӧHt�L�"�mxx��q�m�����ߢ���j�9sf��icK�ǎ+8)����F�������?��;�-[v>77W�����g�v�x��EQQѠ����z�J�ǐ������p"��9)�����_]�3fH�_�~�سgϚ�S���>�:- 'pɒ%�\�Rg�J����H��FFFF+A�0���о�}���ȑ#A�c�E�����R�|&p�ђ
�v�L�e�������e����Ž
�ɓ'e�6���
,%%��~�/_6ݏ
���G�n������נ�"?�a�>�
C�������bt�*�c�C.�4i�E���[�|��իEII�d�رc�.�gY�n�'??�* �[�?^�ť5�(,c?��J���@�j6��k(�ܹs�J���ƍ�ki8����T�Uz �WUU%EEE}a��O��@�|�TߩT��Uׇ�"�Z\q�ڵo�o߾�-[�t3
��v�F�+�����ͻ�=�hGAa���U�V�6O��P@����/[
�B�(D�S�T�}�'��;��m֬Y<�6�fϞ������>x>��#�tX��v��h�� ��s�Q)��y�w׮]�G�޽{��_UY*ĐP�F�w|�U�G|��@�R�>?�Q����&�UB #�|G<��H��B_֫�۷�5X>�0a �����!�˖�����VJ�P>Ko�9n�С���3�%��W֬�s"�Lҋ>�9�J�������&aI�f���t�V�"�n��D��3��n�����J	J)�5y����Q�M�:�1���D��8��ʑ���@sp�ѣGK�����4�;�B)��lU��2��=��	���	Y��f��Q��@Kcill�FaT���2�T����B�Æ[z�ȕ�6�6�by�Ȗ�P¨�
�p2,Pưj�8��8�1�;@�o6<]Fg
��iĔC-=����h<6lBm���WY�Q�w.��ssk��Y�vc=��
�#�V�g!�����}J !�	
1����P�����(-7��0�1Ɯ�qX[�,�%�N�t��R���,���Sa4�b����w����'(������N��ƌ�a�g��T]�*V���L&q�b%e*�c�̻����TN�3���cdRWHii�T
������N	�ֆë,�U>T�6<���ca�ň��>�MX��k@&�8`8��555��Uk;�1A��4)T�P�)�k��4�݀j�ݰY	4Hdeeɤ�
b����ʔ��2R=+��r)Z���f����x1۶m2�he��ׯ_��X��}���LPj/
6��P�f���~
�8W_�c@�WH��̒/����7o�,C
!�IOO����	ci��n+��P���UکS����Ƣ���ۅ�����Ł���0	�6m���K<ً$�ݵk��R���JVc�Q�ԯ[���
��v��������G����ھ��bYYY�5��]�����͛��!�?"@�2c]�$�PE��D�P�
�En�ym��N�/z�������35��T��������s���S4�l���f��r�Y��W̓^&��B(ߏB�`����G?�%��_����Ez)|��M�J�4��D��.����ŧ.�B8�6//�h��4�ҡ���R��C��q�j��J����5�G��ّ�s654o��ish��J�YW�^m3f�^�c:�����"L:}�Y�_���9O��z4d�2�O����O ��'\3��x���x�-�?��0߁Q�f��$��� �JJJ�V?
���wϕ+WDo�U�Y��B�;�xIxK��@αB���ǿZ���+^?O�;yF�'��\��u��?���Sxh���)	t]ߛ�_�'�S��E4    IEND�B`�PK   ��{X����?  [G  /   images/55b8074f-3515-417a-bf4d-91f9a1b9fc8e.png�w\�]�/����B�&   54�(��- ����R)�A��N�	(J��JH� !�@Ȇ��v������߽w���>O��9s�̙�Μ��D_���f-�G���'��;K�΄ɡ]�?״�c`�;~��BڹG��������������:1��yy�9<{�$��뒵����p�A��}���ՙ�l���e�nc�S�Q��N��~Z�M�,N����>,��ہ7�n��Iӛd��b�>�[��ዎ�տ{/��3���J���s��]8:=w����]�02Q�+�Ȅ*�(�(㼣��2s��A6@xF\���o�~	��i������j'/��8���pR�N9���x|�q��~������������|�_���og�Q�_X�e����ր��<s�A����S:[Q����b��O��
X��T�6�+���E,0�!���{�j$�J���,'��p gUM�Q��5���fTR�1Lf[C"S��1	��ӌ�;?+��G�����
)�e����y�S2ۡBp�/��di-ep�y�<8=���ʩ?�k�|�����
Jӗ�V6O8O��㧀�!�&��!Ì�!�xly2�"�g��ʿ�B��~��U�����-)�4�p�A��8 ���f�kԅ����,�����}5[$氡���x �eRl��D2��Œc���s�u�2�Ox��M��Dj�4��;�ۈ�F�$���]cl6Uǐ��ŵ�L��_�푇���Nѡ�P�w|s�	��bC��Os��s2���y|�����X���z�|�)��~��۔�+� �
�q�q��dv�ݽ��Ț���v��d����x���k��^�(�O��z���	|{��l&]1��۶������vL��U?ل	3Ԅ�q�_�O�p����}GLZ��
�9&w�FM�h��������T��M�vX�Q�����#ӸF��v�?������2����O�Jo�+b�//�Y�{�h~��vgjkA�)�g��Δ4���x~jF�������k�OˍO��v�oH�mh���ϧ�l�XF0nw�������n6�=���d�4���	�;�r��Zc;��tMT'g�V��� ���:y�h��cd��ëɃ8v��G��Jv3���]�0�Z��:Py>��7�`�#90�CB����E�F`t��/�+!듪�Zr`���F\�򹪙��y �2�� ��SX�!�N�i��F�V%pZ���l�����&z�T�:�$�TlJ���|#{F���Ư0����k޽g�oX~���&?�7��_�H���_�cY7
���������֖���$���
�A�bB��XN�L��ڂ"1��^Y���z,�}lT�ڝLS���{q����-�K��@�p� :�*��X饸�����X�k: ��j���!�z+��qT�q�Y�߯W�6�U�oi:����v＼������ �&�?�v�k2g�OT�oj�+ *�#B�>Dr(/��]���N��ʶ%�/s*��C�D6�n7_d[aD|��8+�RD\�:�|�(�O�b00��N�K2�W/��5U���LݮKF4��X��o<꯺OW7� �����ڶ�I�W�T�5�<��S�����T}7��Gu(�^�������(ڨ�[���ap�|�9�h�$�-�0D_�J.����\��T�Rs?�!@q8GG�܌�4Ý��(lـNPx�v;kwXm-���k"�N7<�y�(
h��;�[����n��#���A���8�{E��/�� �m ��\`C�<>�E�|7���n��@�NU�n6rEJ��d���A�HY�m�4��fhjI�H�_�5���	G�;Ym˿����X?��6�3������bY������������'.�V�6O�ҥ=�}�^�JH�xᢩ��`���;�/r�~:} �SȀ�ϓ����Dz`Kv��䉈5� ��1������h�qs�Gk��L1c��HZ��g���y^v�Қ���hW�I�"��|0}�i�&D7�f���mcF��
Ǎ�Ѧ����_R�����_�O��􁦁�І�n*o��V��1�6F�-Z���|-(��[D���L�h�۞4��_�e�&�-�
,/}�_�юTk�S�V���ϟ?yHR�碣\>��ʛ�R �9�q���u��+���&� ]����5窟=|+;��O��-�b��^\����/'P3�����ܫ%��gBl�Q[����f'P�[R����ۃ8�d�����tl0O�1<�X"��Ү�䒭�&�\�A�7����T!��k�tu}��bs��X$�(\t1�n���E�s?)(/NV�9+�B}-~�'�ѽOr�]&U[���#�7Ԓml>^�-�1R�l\�_�G� &���m�ņ�������������R���E_i�0z��t�=
�j��.��m���@C��>?\թMĭw	(.Uy�M�W#������&ؾ櫧l���e����T���bU�l��q3�}�������3=8���L�z�����7�����/}5-h�����R�i7��dQ�`��~�C������������)
෭x���!���V����T�ƶև]�/�c���cԏ%�W��!d�,������`P��֬�#Z�Y*�]>33�B_��o,���5��v6ڸ���p��顅hҧ��a�h��ĩx�Rn�ê�|:�*�'�]
|ҿ���#e�Β����9�����V��s���k)c�����`$��M���Ud��ԇ����e�93�m^I�S(i��AS�V��������Lp3�����.���K�6B���ݹ���M�D���
�'��LՀk��7Am2�3�Y���f~�����{\?��@;���ίL��q��b�/��
/y�Z}h_} l'�	�u���Jxrg��<,yp-Çu�
��9J�!�����8��R��l)(++�]�Tt9@�1+ta+#������ M��__37J*,5�pm!W�� ��M�O���٩qppBm��2�������5|��a�2Q���.��/Ʈ��8��U-��̓��Uy�l7o5�j#y{�
�׽�]8C[��B}6踟mN%�"�����f�8A�S�#��iQ��0V�aק9�jD`5�ȯW� ۜ��,�F\�r����t$0�1c�dKf��g�B�߾$��o������T�<�G{ş��`���!��|;\�������-Z�?�m����`H~�`}�7�nz�`C�C�޾�U����7.1aww�H�~� �]\I]"V`j��5�f
U7I(��q�ߗ���|ىI`=��X��7]FcD�pP�6`f�4��β��ڊ|�j�g��]�хe&�Ω���6(�w$�I�W`��g�T��]�
c�3ۭo��߻��E��GTt�x�hyi��#c��f%�;o9�2E��GO�^�^��Q����h�e�YSUvu��d�������'W�)m*T���
f�\�<�?1�]ï��곺m��R���ߑ���"����T\�vk�Ό�L}N҄��Ϛ�5W�\*���g��Ъ�P��ofsp�K���b��~ŋ��B�Al���x�H&���?̹����zv#�as+�����Xl��Ƞ�L�fl���	&f����;����_m����+j�U\��z.r���냊t{��Q�ūJZ��l�2ޙ{�*K0��N��c�o2�F������î�����}�ΌR��ښ�>���O~��i�F-u��d��s;_�i�*7����0m�W�(3-�vP!R}�:�'��];�D����|�I�*Iq�K��W�E�!?��6��v�FZ��m,��E�2�[���8H��&�!��}O���S+��W��G�S\����U��VHi����_��X� p7�(6ല.�2�m������4�������1�K^���ʒVf~y�I�"u ��D=\���.��+%� Ga;�^��r*��Ҿ�'���s���u�oc�J�J�ugO���Ě�J�����np+�oDs���lw��+��PK�+�C�8���hx�� g��d�)�{pD��_Ƙ�0'�)�z��R�J�%%{�|e+8���6ǿ�m��d��=���/����L���> [���N�!�C/������/ӫ�=��36�h�r���w��ǽ���s�s��|Br7>�u�B�!.)�	�ڟ�P�P;����Q�n6�{�(x��a< �-��W���}�3\�۫���H1��|�̚eN
�	Z�m��'v6g��K`�3��l���/q���ޟ�����/4'�䱥��E����d���N�a��hs�L��U�H��p�ĤQ�vx������Z��^�ÂF���~�]�RLa�_4�!�埣'��?��sO�)�4,�����ܪR�h	+��o���z5��{DG��0�[�vG_��7j[�E�����0�V�������L�Ay�����ư��c7K�&�OHg-�}�}i����-�v�[Y��Q�e5bt��e���6n�3����`�ӫ2�����ޡ���5�T���Ǆv���%?Un5i��҂��3��x��x��˞(-��Պb5���q��Al�O~�ٟ�g����^~��!�3*��n���z�ȯm�P��O��}�l�x�뾯�[�5m��V��Uq6P.9:�/�w�3R*S��ll� 9���芆�ш����Ko���C
���`E���g������i��è�X�!����TN�op{2W-�ln%_Y�<�.6�81/�����r�W[OI'.�?
?���`ri]@*��Tf޷��vf�cq:��2�N%��r�O/`�s`~��C����(�BvS�1�k�3҉����V4����n�96}�y��#h��<���`m�MO������1�|n���G�4Լ���/5��-�V�%g�p�(���q�����}�3��^����*Ї���vcqu��7ω�s���^՟}�o$K���o��˖��y�����4tFP���A\5a�o�>���K�h`�z%���l�=f ��|�f�l��P��v��Q�P�:
�t�xL���&&SI��C��f�ܛ�g�]ޘ������r8�`%/���,��?�@�ݪ)�U�@<"ou�����|�Հ9c�G��L�ʒ��{�UA3�U%��9����E�d������;q���[�Q����")B)�P����[����<3������}Ve���H��+���m�=�Cr��Q����t�Z1�����5	S��2�u�R����]5���<��l.<(���ؙ�r􃇯j��'�s�^���f���5����΃������5r����y�6�yo	.��O�o����' vEﮍ A�I�|f�+���L�I�ir�P����/�cu��5��<�զ_�8+%;��k�8m�j.��ԇs�%gDzF�v��}�����~U�.U���w`�b�MJ���9��#"�j|VsC?j�'Oph��#d��OZ�k��~���"F�z�I��nO�Cay}� eS������w���܋�af�h����mr�^�k^�͡ߣ'�ȵ���E��%+r�~ߘ�GM��t�E�CX�̫�s73	�G-.N2Đ���f]L�Gb�J��7A�K{�3��ށ6V��_�=Z=�"6��Y����y��ޓ@"����de\V:����	F]�V?��VVm�==�����χɅ�x� r��mqō�p���g?��7��f���x�W@E��4�QRIW��<d��s��������sf.'\�m<�I`X���d�7h�u�ݲ�Џ��7mϵ���d�tD�y��B@�� ��UB���̪��x��鮴M̧�+5-?�WӰZ���z�/^+ ��'�=Ό��~��wk0C�Rׇ��]%����a��/̎6}v�}��
�r5 �Lp���;t\���1�V�����)V�����:�B�fS��G�� ���1��\1�gZ�^�X�i��.D���۰���d{s��7��3���O�S<�4�|I��(�NiwV�N�5\�ڹA�{έ���x+����p�?�0�,P��ă��Wv�'2��rY���&�#��!ئ����7�-����R��Y7�m�!U����Bx��H[��M"�E�X�6��v4�vd��+J__O�`]�ycf[9���<XM��GӰ0�#���B�_A-�EE5��������K����#�P��qo��/X�]��f3��Y0;�r#DG��B�8в��� ��n=�e`�7�}�����8��L#[r�Y�y"V?��'��Ȓ�� Ő)�L��&��#�p�*�\�<	-s��z�lN#����]���
���Dч��Dpn�О��N晧`Օ��>|ժ�0^�T�
�Re����	;��I��Tl&�9���KQ�!��.�@I3&ؖ�Z�6�MÍgexq3h�MI�y��Y���u�?oc^k����X��8���˝�m����Y!�fW����>Iv�< Oé%K�_����*��5k��ޗ|�TQ@9MAa'f(������O�_FuY��i؋�'l��f9/�M-��E|�) %0����7�%�^&{��#Ԧ�"��*\?~��0{D��Ʊ�+T��J�]n^/P����������a	��;2��A?@sqg�w}���E\΃�tb�q3��ң��� �W�_�K�	�)v���g�<�O��kX��ޞ{��H���lK)!�A1`΃��%�~b��a�r(�#{d�A��vNw=>	iJY��6[r��0y�Z��36��� �0�r�K`�����n��ER���j�^�p�<��0�6�N|�y��tE/E���,-}����i���N�e߅�^��7��}�2Jp�mM�[��\B-�< ؘᩫ�%ѹ0��uދ�W~���f�n��NDǭWy���2wGl� �U,��ݍ��S�"���P��E���cp�����23(�p�j�꟦�ʹrɛL��rƭ���-ȦR!���[H��t����~�ăS] �`�@��[�-�k�B��.��X��&�x񸽃`[��{e|m@��p��vaO1�Q��h�w)0��{ҕ�N@g��pY_�{�qY���S�����hn\E�h}�>��;��˖U�/^���M���9N��&�O��:�/�N�L׵�4V����|��\㬂��:h'����C��hxcvT�ߋ���
��2�D�&��,�w&Q�Fv���-�V�a�����;�0�?��X�ͫ�^$'Q!��K�ׯ����9lM�LzdI(3G�dv�V�P��̝X�K�so�/��!l�N�5����"h�9����&2����JNS��Y!K�����r���?Ձ<�>��H�����piA��k�9��i����>����e^6z"]�,�|�o��n (��ڏ�?�=��Ӳ���|eU���[�ᴙ��@9����܅��'G�`w�����Q-�\D�{�m���ْk�5]���#X�ԍKϠ� O�y�vl�R��3�>k�u~�>�%w)��k��~���:��UϖW��\><��1����2,�fWR��Ө�����#�s�� /��*ʯ�x���hsa�F�l�(Hĥ����H���?��s��DKߪ�a�W�[툣�����%Z�,|R	�����ƚ}�(������a��i�JL'�<�G�Db�k�~W�Ί���e��۾�زQ�0WȻe~)D5�+˰�Gx�E]�,4���b�˟`r�����g�b)J����|ޛ8�%s�ecY��φ�\��Y%r�>�ݯXyZ����7�n,�6�ᕐ���������ReE-	%f��ok�f}�V'��M�j�M!{c�J���Wj��rKh�����߬�`�����"j�/?��9���韺k�k
�<��/��ݡ��[~��M_#��K?Xy��X��D|����.����>@����aB��9�E�Yx"kK�t�P�#oJq ��'�<�72O[ ��};�����Ȁ��o׬��ՙ���F��?��u�P-��ǟ�0����U���r�����)0$����9ք���-���5�4Y=�F��p���7
`�j��4Vz�e|��m�.�U|�ʺ��i�M�)�H�{O�"�]F�9�˺�,��:�%T,�;���:�`�p++��#ĬC�%�P�?�L��q���7�, >��?KɵwJF�G�������Fy�G*7����=�����粌�l���G����T��sF��3�����W���a �W���|!�)�֍�g7��#8�ۖ���'����Yo�<=}�>���$��T_n�'�憠;������~~���+e19-�?X�a�'�/�W����������	��-Fv�ۋ\ъU@��g�5'���U��2L*y��Q��fk=�R�n�VKadH��$��<�X�K�^(^�{TN�l�O�Yo�i(�l�=[ƭJ1��/����A�<k��!���wg�Z\� W�[�=2����ӓ��3������%.z�xx��w/J�K����9��Hמ��/+��	T��,�Ҿ�-I�{��e��ͨ�L�znB�W�(��ʺ����<@X)�^���ʉ�]̹���x��.�L��X�LtQ�R��������3�u�MI5iX/��uZ��V��6��u�U��s�$4�e�$��`p�����9��\��J��DQ����0)?(�	�dw؎a�<pU=��?�b|�V
�37�djߟs`|��#鞷#iwa;���ndG�P���z���x���zuV�BT�bu�T'�g�@L��$j'�"/����X`�L���)>�5{��Rv�#j;�ztΡ*��b(F���K��b%=.��T��Z�L���S�b����w:[/�w����d�6e:�׉����R�B�9��<IA����~�AgA�:¯8�/<�͉T�!]�hz���^�8L#ll�m�§+~�(,�:`�.>��@�\R��U�V�O|�-�y�d�=)�B�.q�ȹ���[�A���H��Rҽ;@�q|� ����n��x���� n�Xk�_�-��u킝��N�A�rw�\ �/��敏_u��e7#}`)���-+����@������$#�ԕ��,<�����'Tߕw���u��k:���}�����\�}8�0Ll�@�"�a���a�1�����嫧���&����u���mI4���G�Sˬ�鏓~y��"r���=|ex��������?>|n�ݤ
�OwM�lb��'��x1�.�;Uѐy{�	m�bC��S�-3\H����TιD�}/:�+�/���T�WvEڞ&�����Ν�e$2|�����M���t���ʺXC�r���.�\���<SVaɇ��YO�,˙D�*��}��q%'l�ږhR�F�80�a���q*s�t�G�yٍ�$��N%�Pw����A��7�����z`H�QJ|�ك�oSWiC�Iw0�-O��L<<�z/����3�}��hAJ��
\_ܮ33�1"��!Z�a�T���;����0d�ZY�����3�.s��G�(���ط��j�m���:s�P�MG����d&p:�u��WedM���f簎����U��裍�����b}f�}s�m�ٷx݈������5ՙ&�yL8M#���8�������Sq�8�P��w^,ߕk�XM�I�tW��
K�as�����y��QG
��Nt��pȤ7ޖy��Q�l%Q�l�Ÿ�=E]X��sfx�k#l�݈,�p�;m�@��KN�0�2�Pl�U��h	��������\��x�6s�H��M|���r��0S ��B�����Yٸ�d�ct�<����gK�z�����1��H�aK=�����"�����L�@^��v�ZZc�(��MM�j=�0�mÝx�>���� r����K��^V�u^� H ��J�r��
���W�����7�x����P��5�[����7f���#W�vqia�ɡ-R�Q6����#���Ѝ۝�M�w�b{�%���v�f�k�dq��[x����׈J�e�����>##&�����"k�ŵ�*OU�}�P�lcX�!'��Pw�B��G=FK��xCh�2�m��N	��T��b��?�-g�R#�-$�l<`Pz�d��<�W��Fܸ�'�#+e�6�-i$d�[�<	�w�sA���2����|, �ѷ����
1L�s���-o���0��	�^8�TƆ���[KQ�-n/_}"FHGĄ�I�-}x�՟���	N�f)6I�	::"�=�j��;���t�:h�\J��3��\PJ�mSU���O{�z
d�T��C�+'-NZ������:��r�Dy�H5���x��M�{Љ�D���Ͻ�5g�>~,�\���$��%�IO�P�sw��b曲���Q���c��PE��p�@pel�#�&D�1:��*���a�wQ��Lm�sH������Z�!����X{�M�JngE�����`*,�8����yw�c�VrC���;���bE9X��#i̴�x�?,C��	�$X;L�~0��RL��m����=�c�J�	^}�����@�� ]f���@s���o����Q�Ys��V.���R���������]x�ω�;�B�R,\�H��|��}ʱ�q�>D/܂�u�1GXJ�4�"��d�*�~=�Q`C;a�z��7���~0..[�v�ƻ_�P�PRR�sK�j�M����	�M���^[�J�) A��������I%Ay�M#~��Y�pIY�p:j�̗�<׻����#�B�W�^�������ٜ�~�zG^E��ad1"��O6�cv�L��ަ��"Y!-�WT������+4��%|쾘�}�wu���]��D&���V����1fDǷS�{6�����b��J.�����1������nQ��y ز�J���`�bЍ��?�;�>1r'3�i�	�4����Q�Mw?G��7)�)��@B�+EEyT�%K��D]�,)j��%Z,D��*��\k>]�� G�6��1�TČ#	��f<1���5+)�V]]�on�(o.�QQb]��J_gק_3��|�8�Ɇq���$�?Q��4�Q)�}��(���=��^j���]0�IY>���}D�K��b��%4���M���|4�V�~t�̾yh?�����:�|e�q�z��R��e���(imi�������Z<y��	�%���n�Rk�z��C���r�
:̵~��yz�c�gӺ|�ϙ��
�2㟐!�����X����%�ѝ���:���6{7��o�ם�oU$�yƚ�e��Q�r�N���9%�&�@y�kI߃F����R�_A�Ɲ^Y.���;X�P��s�_c�]k���EU��!'�u��م �I2�T�&i��TWJ���X�Q}��o=<�:�i��8�+Ԕ�����"Q��Б�z�׻��﫿���Q{��t���:Z�ʤ\��r�����^x=�.'���D�ޅI�+��8@���ٺ�^m�b�ӝް�%�V��]�^�s����Z���g��ßN@/��� ������W��؅�c4�!p�.���fk���UH=�=����y��jM�ȹ�::{���r+��r�����IIz�M�Ka��|��FP��D�g���ЎMn&LՃ�����o�\R��zY���c��GvI|D�.d_KV:��]����g�	�ʱ�
;��e\�s�8�<sΖ����#)%8H��U�~Okb��9�'С���1E�Iĩ����^0j�_F���m�=��z�yrMe]��s��1����SW�a�
@x�U{'�������28OIbd.�;��G:�PчJ��,'p�5'�����.�6p����̠y&�� ���lO]��C9��Ek����{�H2�:�]>�pj*�"�[�r!�#��0�=�9����9ntͷ�}[7��m�8�3�k��c�=�_r�Au�{�~'S&��WLP,렷�d?�L��9���$�Z�eA������5'��pt��s��u�Cd)�C{��DH4}ھ�gHʕї�H�{SE��Ʊ�����WL�*��ϼOC�X�����pW�pl���b'�厌Kt����:��O�v-�������?�Pj����a�6�dKM4b�@��ӿ����b�|@���V�NqӵD�>�12V#`�;Os�ߦ�zI ��5T}��=;{e������E /�`�jV.>S����(n
���_�<%t�=�)]_�)������w�p�ԇ�{+�~5��M�vh?��l��/�ŋbh�5R�?!>X>'��[�v^�����u%z���;�,�Lu0�g�@�;~�ϩ凄��&�w�te��r9��z{�*I*{����!bν]@�(招�����a8��[�Sp�Q�d�=��o��`>������e>y;N�z�R3q>|�����~)�Y!q��n����E�,(���&;j� ��~��E���m2����5�|�&M���+r �W���]�J�)��=^I��8l]���˺����ѡP���1�3uD�$�KL�O���$wd
q*����1���ꆈ��������(�p�RR?�!�F��G������('��O�$ߒZu��{�6�iY�����6R
��ft�I_�� �>�mi��Ԙ�����Eu�A����ȋ!.�[��N�W#�#�et�?I:p��T��Ӿ 8�Co�i��6�}-�O�?gf�SRBOo?��5���6��7ԍ�I� ��}���;WM��D%L��LU�8��U�
��<Ȍ�T�^v��(��#=o�*�-���S�"^IY �1�Ig�
�Y^>�}�в>`{�O� I�&�t^%+�G�~×.�P}a\�r�ے�\wmc ��yN���z)�n=�&2/3�,�����Ɏ��ر�G)}�;�����V:!E��}����u��e��hF�t�9�g��*����>O᧥��k�]{Y���b� Kh��A��v���Ğ
~�:�ړ��:*�%�0����gRG�+u$��W��VT�[-�
:lD�=�>_r��Y����Y<IR}�Ӵ�Ra�e:��<Q��� ��ZN�}=�}҅�	��0K���Ug親8x6h��3���?�W�kV���	���Q���W�S�,��Va#�L�Ie�@�'�3�D�&;�;{7�޸G���~�Ho�_���q2q����K�v��-�*|y����E�f�1d�������^y��Uf���,���/q_����d?���+�����
0�F:�[�O��oso�����>)���nڹ��@y~��<i%�+��4�U��(��q��\�U_ ;_6ߋ�\��E�6?��Xg���͠A7�$i�ޞ �ZA!v3���||օǚ�WH8pJAn	}�z=�tX�{�q��TY^Y).��<�'I�6��z�E[H��M^;I�7W����yKZ*_��@8�+�����7W�,kj��]�B^�,�o�s�4�K��3%ջ�:��.���X�Sv��6}��?����#�-�g���K���/Y_��}��PVZ*LS����>��z�r�۷��Z��o�wہMj̍����TV|FXN��E��ӥ?8�j{Ŧ]���C7�K]����N_N�P~I8�K����K�R���/���O��e.Հ�SWK찥C��b�ɽ����tqth�.�i�o6`[��~8�ߓ��q0�'$�������̗���
/��i���$�-8�\� w�_�����奡	��Ѯx�?�.}g+l�@�=�=p����ZX��V���Yb$=2ݩ���^�dT,�ɼ�ۜQ�]�<^�{�.�q���o˵T�v9�����)3���i�Jz���3ww�����l�%����iz=w2G���ʟs�j���x}!�{��h�]�	�%%���FFF��=�<V�C��?'+DR�9�؞~\��*�����
"��/(�H1���&{�&��0=���W5=�59c�ʮ���]z�m�L�˳&�}^�����<Yd]������E[��Lt�L��z"`�r�<���>�zeU��Q (!�f	ڢk�.K-x)�T~��8�fo�^�e�?6�M��R+1�c+Tcb;�Α�g����E��������⧘���� �*r�dr`@�:+�[�ǖ�#s;��p��<L�	9�me���_�q���E~�������#���U�<����,~k���R��;����S&�Τ��w�K��4��޽̓���*������@@��w���q��E,�����O�5��co�5$S/n�Фy�/'8^�-T�/�N�]����r�fl����G��+|4w�s���u�a��y�+$���M�pw�LF�����GY�Y��c���C�'�������ր��%]|||&Mhd�鶡�@.tn!Z�%[�o���h?��/w���hO�G�xڲƾ��V��i^�s<R}kC�Ջ��F[k�^�I"qO�Ύ�pb%lt�")����V���N*��C0��uJGo�[�C�y�-U�ևYbC���R�<�q倅'�E��,�Vb�Ј�΅��uI��f�!��8�w��;ſ1�lY	�=C���2�RÓYh\����6*���>�LG���14麇Pc��Vk'�y7�JI��v�C�H�+���/��S�xg��2��dq��,O�H��d��(V���7شN��oF�L����r�R)�:)���1��܈2f�A�=�(e|�#���$�Z������M��w�A7��9��#�K� !�o�A�=�f�|�+6��\�jI/=���aC�#�R�ԅf�>C-�x2X`���]�)�x&f�c��A�f��P�aF����%�G���d2���Aƕ� .�9���0��0�[��O�W8��8�Qk�u�H�ċK�b'��~�x�V	d��	�8��O�%����CŻ�����Zu��?&��X9:Ԫ�&�E	���V}뾉+,k	�by��u�c(��6���N�mI�-���ILYX�!h���e�������c�y��u����_���!�0ic�B4�I�Ξ	~�a�X=[.�8��nO!�U�I�r��[�b	���Ѷ���_Ðȧ�<7����k��V�s���l���W�Į6%vYu�FB6%=� P��cs�qc�ю�ߣ��ƌ�c� 	;c�+�[�X�E��;ӑձ~bw@���~�u4�r���[�z�ue:������z�<)fM���-���d���H���CCk������' �z���B�r��jC!]]G�O�h�*λ���5/�7*S������#���|�u����Z�{=��o#@b�V���>�
"���mg�;�$�]�ײ�����:9�B։�n"DۺS,��Y��^�����G.���"�jW��r��V�L��@0���HD���(�(R�̃�k��ŽF2��7��F�!���^+r�эM.�c���Ճ8chU
�&���7!����+%:�Đж�@\��e���B�ʽ��l'��D��;F؄"���M�o��"�B`7>Z8E+]9(�b�ËE��f#E����5\2�x�V1����P�H/�,E�^r@B��̆���q�=��h=�J��[���Uce�5+X�Ɏ�%��
��Tyܖ��9�'5�����k/�8��L���e��W��9P=�픅��o�h=G�݅`����v^�l��Ţ�.&�̈́��&��f+4A"w����daU4�Fv'�"����d�_K���[rPȴ����~�g��7�Q{��2���k2��5�(@s�ܠ(4З�O�a?N^���k.��#"��g!cr�����?��x�{���JӶ���M��Z�����+H=���hs����|Uނ ��d]�(X���Ϧ�;�O<V"n��}^`_USEdFh���Wj�Y4���5H�K/8N2�{��)�߯��$�4�4�0th�4��n6p`�K)��-�R����Hԓ�q�ՙI�����c�G��^�/PK   ���X�?HU!  B#  /   images/585092fd-6de4-462f-8499-92296fb2c536.png�U�S��]:��n���	i�F�;�F:�����n���n�x����	�;s�ܹ����=s�<��@lJl   TT���� $lL��m�����EA� ���o#��hB�]R���u�~�t�0q� xxx��8ڹ��|����l�y*A	 0�+ʂ5=�N�<5g��=k�K��"3c�����s�zhj>����v8�*����U�]635����D2a���Dc������M�P~��"z3����l�Μ�ws�+<����1v��2nh���0�*�� �dz�̗.�`;7)�G�fK{�"j�R��6G��e��o���<��Z��o5І�h��+u�8oi~�'�f;- C9p�]t���F�,��0^M1��D�K��7T��*��F&���Jb��{.����a���"�P�R�9)��H��G��3qx�N��
����=��Sp�IP���=YQ#��Q-��\F�A� /R}cЩs�@} 1���H%��4�k��(6K
w�Uxt��c��[?2
��Gh 6P_�-���(�QXA1��+6o����ws��p�&E�{�Y�X��"�UPӊr�K��=1��8��K�K o��H�hV����[9�p~S��}wuZC�p=3��GPZ�d��-��jn7��~�ʸ���O�֜�����3iZ]2nT�p�'/��g�}�iU*�k�u��V��gOaG���:p�r�N�@��^\��	^������N��ś���4��Q���S��g�S4O_��&�\k����ീ�A촱4��N��u3k&lE�&K��q!� C؁HsCY��ۆ�@�[<�I����|�h5�@w��6�:<��#�w�\�ն�iI�m��G������,�}�f�ԁq�cc}�zu���'�4�6@[�KW���<��T����4.IōˍY�*��1�ف�+���R	^��>�]Ư�;W��d���tV5��C�xłyx�^hE�윽���d���7��7�S�+tP2�]��1��E�9��j����60��Aʗ}�e��3�vi#�k�cNv���� M�U����D�@E���y�̴o�U�;�]�t��n(-�"�B�}�2v?e���}�;�{��'��{�A�/7J�3�f�#��{2���t7�0����-��'@~z������
 K[���ϗYSIܯ�K�>���@ �p�^��z�k�w}�}���f�,��sT�yzU͑6�3s�7G@k��1u���ˀ�k7��q�������������>տ^���� ݔƥC��,U:V��3]�u�������&C��j!���W�>ȹ���/be\~Ii
�l+�����`$E����Χ�"����O*������|䢤W����'mo����
��glFE��_$�)�xK�EC�~H"/לiVcƁ.��4��tFNX�/��Z�3���Tlڶ��đ�Q�"F�VV��ե<_Z��������X�>��ADr�_��-��2�M��[���Y�£����R�"����R����}�$�b�E��x�@#���H>g� B�ӆ�z��F�\��@tR�>��d���9�����8������N�1~��Յ�ly�H*�n(�d5��cؑLG�s3����j=m��� 0��R�ˋT�eM�-֨�B.u&o]��?,��aGYA��i�L�s�x!�5�7�������hpy*-�l�_�FӹaQB��s��c��ٍ��4?��\�uO��`�j�!�����|*����P�嵙�1�@m�º�t�:���g(�<g�3�=��u&?�[GG �ڗ���#�ڐ4�Я)ٯ.���wޅ����0����(-�A����yC�>[}5||���[�
}	~�6T�J���9��x�x�4DE�|��_.�1�.��l�6�Gtj��;o}B��@�����̛��/R��J�q
!3�j0���[@2���}8Cv��\�MV�iM�(�L���� �G/�~S�߳����������~"���
������ߋ5�yW�O�c�2|*��[���3j.-��ބ�"���rmʅ��m����߈dd��$NQP���f�546	{���|wRZ�I)/��Pάk$�3�6����~�RfU������u�ס��R��tT�6�u��S#����zd��y�w^�Y��E�'�����H`��i�1�"+�ˍW����	��W��0r䳒s~�tC��5�n�kZ:f-��j�7��g�q����7��#M|�<����
�梕ѭ����+�E}#
�̸sૃQ�z�� Q[o�伿��:!�ޗ�qꏳL���XY��p;~��~���ΩEMBD�sw�M�!-�j8�Y��dT��k���4	����c�*[��P�4�4�.����
�o���� ����x��t��������ye�o+w��T�g��}c�;�#<�H�<geζ�����_S��R��5pVSP��{���p��7�n��P��<)�ͷH:��uj�RAҦ�(�����ݳ��/eB=�g=v�	�U���62#]75Gd��nt|l��s+��hfn�ɥ�M�N�Om�"�aTF�'?֖旱.��|H"�ǚ����ϛ�>lس�r��L���޷7	!�`US=�>4�煖W�FNú��(q�asǟ�Tc��6P����Ie���1�S"��T.���n7u!�f4����os{kW����/w*�����.��%&�b>�p%�ݾ�%ߌ���W�'����q���O�Qf�B��!n8�sn
�~j~���|7�VU�Wj;CH��99��v��\QA���o�;�S�lj�٪V��Wf4��H2�8��د38�T����ėh#�f[����M@�E�'4�Yu޹�������e��7�e�ٞ�2v�+���?=��9)��Q�#�S=Bxo�k�0֔��2��l�M'}��B�r_�f��{�7~�W����<|KD��-C�4��Uʼ�jHa�
m����ث8��N\����ZS���Vڋ��G���瞾��l��zn����'��l;�W�m�K8G	���[��?�c>H���J0�c�����;�?��w�6g��2��(�1AQ���M�y���[�d��T@�i�-����X[X�B���f�0G�k�d�_��7w���1F<�l]�>�^��M�	��q����H�KzmY�82�#�s廛��E>.&�۳�ǥ�g0c&,h���6u*����U!��2J�|^Q����9:gr�x����]-�*o�F�̱�`��E�@�Jho1N�2[�^S���Zf�:?�t���T�Řl!\X�����
�0hP�"�w{ɭ��RiDc ;a8Ir���f�[��}�o"P�'��OG&$~��4��|nj�2��oǺ��Ye��!�<?��KY�:5�+f
���ɡ�8��\����L�����/
G�C��Բ�9%vJ������X������E���7VR/A*��sBN`L�p9#�(�9���c�J 9�O����FOY��a��k�IƘ�����BpBSLI�*׷�G&��gL�a��J� .�rǥ�6�.v�_mO{拃��~_�,�a��y6��@��4m�\6���B_�	L�𣖏���g�֜疸�TüO}�>�㇁���������>��	o<ƍ�������>�x3���H��Z;�)x��t���v��h䏲�Ws��ѣM�JgBSW׻/{=�6Y�/}�G�a�|Tၸ[3��9ހD�)l��?M�7�\ա��6���]fq�;�|�0@	�/L�IZS^|�a%��Vz�����9i���G���﷞�;5o��.p����7�X`GD`t>�-�Y���0��o���h�p3��r��;z�q�����B���^�����`�vH�%�%ͭv(x��X}�c;����}`����H��yL>0�`��m���[0g��W�� )Fr�Sf�$m[Kx��z�	�۫�G%�R�O��
J��+��F�]v4�9���;I����L���8��ҍ���wN)i1j���c�T&�M"l�"��L7�7���)=\� ����z�g�a��L*t�jB�g'�:2���������2Оt�raȧR��y����8��YP�Oh���a$6�!8n����,?��C'���.�M��#����nj� �~��K�nA�;�k�u�/@G�]S(�<k�lZ��Go��Ϊ��\c�e%�d��k�1i�"�5� ��=��t?���@��ƕ�8v���wE�Y������h*����r:Ɯ?�ms����l�Rx���~���o����~�F	�cں�?�Q�U
!t�����mEE�5qs��u���2�Y���-IJ���<��&�KC�B2���ʀ�]~*IQ�%.�Q>9w+3�@^�L]���`@X4���r�Æ{2�`)��<>nLʾ�Bk0<;���yK����ޘ�J5�A����n������HƗkh�K	�%,�û��Y�K�>�b����T�֓�P� � �ΨR�V���fM�{��;/q,T ���5m��'3��6s�׼o���a�֯b-x�#��}�q�Kv�7i�O��R?@Ӣp���/'e޺"�X��ɏ�����	-�*�p%����A���
�����?��nD��@�\�f�t���7n������XϘ��h_I�ˣ�1!^hf|�VS����.�'+�?߀>��^AP�fg��w��1!蘧qs�����xAp?�Ы�㽋��`z����6�'���f:�8��l@�
˺R��l�@<*���h7�Z���<Xy�{�#���L%�v'S~W��z��T9O���gc���k�U3�@�#���U�z����WAV����S��om�:Gx����U���xEf��b�J��:��,�D���������_��a��N�(����ο^^2l����j]�������#��Z,��^t�x��&x����%�A�9W�"�{~v}����t.�����H��$�h[o_#�fá�<�,��X?hr�x�IȮPJ�n�w�����d�&�(x��L�����K��^�BQ��lc-$����mog��v��>F���}�|�S}g(n�y,�\e��C}uv�i.u�����~Rm�*��MÀ[�9Va�/��T�ę�M��0�fz�ȁ�����E<��??��3�N�+fk%�5z
?�#f�(�*�����z��'�EH�
�:pơ���3tL-�?� ףg�Y	�h�wq3�wY��Ë�R\�d�{�����c{|���㄂<����/S��Y���f������,��C_�Y���Sm���ay��.cy`�n�͘����!Z*L݌����63�us3ˣ�c ��ݵ�h�~C%�A-�.�&��`Ƀi�U�H�*�~r,��i�'a����ӂ�����k,eFJ�`w�5o+���D|d�ɰ�KP��d�:M�`q��~���H�@K�y��@� �cidf�_�=c��`�b�yJ��-O�8k}��b}x@���Qr�bIi�\P3��,�a�!�_s�����K<����v�y;��j�WU�4 {��}N�b��&�$dL8�[c
������*�ܙ�8�B#F4�F$��*�~ᚾ>�IL��D\��7�6y�lHY�E��C)3%�᝶�nzl��ë&�G�$&Փ�B���'�`l *#��͙G��i�7dij�ߟ36�Fs��e
��xW�<Jj�i�y��꣰`\�H��b$����;�c�V��DRŷ	��\U��ͭ��y�آÚ,x�{��K��R?��E %�GU���:i�@Z�H�������٥�o�r������p��9m84!��9��q�P;���c������q�N���`�<�_m�_-�O�}�w\�N�Z6���ƾ�M��՞�������Dٙ�b/�BW�M�XT�8�y�����8CKі���8�h���T/\T
O�Z�V�L=��x���,��x�v����J%D�����i��[]^,��G�����>z�I1�E����'[�4kq����((fܒk�x�`�9�Ń�7⏑�Z/t1�$W���{�t��s���ܠ�UO�s"i���'�X3���>2�������O��j�#�]!���IhJ�D<]���������I�81��2��6�|q�iǂ<���Nr��;9w�=������8,�X�&p`	��9w\
VG.�8.q�EM�iY���@��q�1m�j߅6�}�	��Q��su��`�w�Q�i�[�l�!fg�>��m���wM$D^��+|>:��˖ޫ��Yߝ.6K�=0č�ө��e���h�s�{���x\��Y���*�f����\r.�
DQy:���[t(5�jM���d$���K� l#5�wǐ!��ɿ��Y��D*��;!��!9�wŲ)��
]�Q	�ֿ�/��q���������!H6���U�o>1��A*CP|�g����)v�J�������~A.-�rE�6.�(����$.���H�)�#t�U��+� �G����_��?���/�~��fO��)|rn~���S�Fo�7���R5��|���:�?N�d��b���g*-J�[�'ʺΝ�V���0��KӠ��K&H�'�������V����!��rC����ڳ˸��|5i�r$KȳA$��r�h�P�-T�'z�g��@�H`�;�<)�E�>��%^�H�6����n�����M���r�\�h}�*��V�4��Q�	����G������AR�M��G!N����v/0�����zy�����Q�!�WNqY
��o�04m�[�9�qQp��o�W�fSB(Ku��#�<'��'ϭ��gB�_0pA�bٝݪW�FX�l��I��N���2�&�?�����0(�P����=]D[�>302lv��̫��<⍌�^¤��q�Z�О���Jі�H�⿷~��[>�U�R lļ�R$y��!*�(ǻa@}Ne��`&<�!�I�ʐ���ć��m����+�&@�E'Hz9b�o&�R���&-�v�hyA��<�}B���Ҥg�(�!�%�jCP!G�jNnnD���ژd���.Π�i�U7L����\[���	.����!�A�{ Q�Y��?m��ak��f�1.00�S��!�sSA��f�%�Np��(�����-<��t�d ��0���	j�$L;j��
�\�p���ڱ�������{#8�x�ˌjN�TnU��f4��u�o�9�uD����F<R��e~�>�Kb���$3���D��x�漹��h��x4��a@������_Fc-�(��7���O h?��~I+6�~��/���h�Y�i��_�A	�������eT�$Ўl�U�3:
U:�P��W�6=��8K�V��7yѰ�*��$C�O�d�J�D-��M�S>EKN�*%Y9*�B絥���*7'n�JI`�CFʄ�w�����	C�:�.WP��1%�3	�[�lC�V��G�;�h�Pd��]4G���P��l4�=@��2����?�#N��µ��F��!_�Sm�4����dY���+w��V�r;�Ovd=X�~ɠd�3(,�WtL�jG|��/�B>�Gi}%聖3�1�T`~�#$���I��a��AN�'���,|bHM�3�-�"_�_4��1|���P��8E����,�@J��X*[)<߁�2���r��B�¼#�a�=�%ە��A�Wߝݷ8�^F7�fz��R�b�M�n-�k�A��\t��_P՜~f�MG'�sg������Rn�7�Ѻ����"��6�5�;(���~A�nԹ�
���s��6ݑ�����Z&� ���c�I�y�?�l����ђA$�͟��9ȧ���f��cPUg��	(u�>#
㏾��	gA̡ɁX΄ZcX.砮���hT~Q�v�z#���ph��'7��Z��Y��Z"��Y���b��p��2�s����hS5/W���G�h
=�=ZY5'���4��3�����WY'�����,Cf����d�:���*���#�W%��W�x�s��_U�I�홗�����1\)�e�Er,s5�r��YH�H�q�1û��@2D�R6���
�6y`jWDA2+9���Kf�L��9l.LU��v.�@�����x����X��񪼗c��`2�(	�N/΁����΃B�,��F9S8m[����Jq[�07w,+��
zE>�M@}����V� K�ZspK�	�щ����M݈�D�-MiuQ�|g�9{ٝ��|�C�o�k�n��Xdy*@��*m�����R�g�1R-Ks���9�d��j=s1�m��x�sms�O�1��[��Te+!�A�PK   ��{X�c^��  �  /   images/817a53b6-1ac7-4961-8971-5b4538e0cf16.png�B�PNG

   IHDR   d   s   n1�w   	pHYs )� )�;d��   tEXtSoftware www.inkscape.org��<  JIDATx��]\�U�����@43\�����
�����̑[��Ie��ܳ4g����L-7KeȺ졌��x	p^.W���z��}��=���s��ʨ�QXX���/����'R��p:s�M�>��ܹS�Oip+�V�۷o7���w���S�R�fef�����?x�@���@\���z����}�:��z�rC�8SS�++�6ttr�Ӣ�֭��x�bj׮9::R�^�i߾}Dj�OM�F���),(���X���k�(.>N���ѡ�ݻw=gϚ�9s��|�]RR�~ZZegg@���ED�<C�;T�����JCC�D:::dhhHfffLF������ٝb2N�A��\�Іf��(6&��RS�b�J:D�biﾽ���+����hݺu�y��}�֭�111���T����|1r�pGW�7����ĒE��M��M����]�6�I	nӺ�a[[۽|��={��0�L[�)5J!���'�#�Q�t��	;g��~~~��z���q:�L1͓���RƒB)))����q��U�#G���ܹ�M�^mӦ�6s�;xv�\�n9�8Ӄ�D[�!5�J��z�n�N���x���G>�ƍ�/(8�099Y��Q�(��ZZZ������B��}���{�� �={��`������=y14$�\\](�A�hguSm= 2�̝C�ƍ��={�_��r����F�ٗ/\#++��I(ؓ�Djkk�����1P�h�O�>mx�ҥ�G��R������������߿D�U�hlBb��
\����ݤ��fy�=�z�uYNN��pt��!�?���I___87n�@IOOO�����`ǂ4BBB�:y���ɓ7XXZ,hаA�-�^�����Q(!������h�z3�f�'M�4�ܹs��5E�C�,(�	o
��i�_��xݤI�;w.-[����&�fY��Q|}�����;v
,�,�5�k�+�m
!�.#=C�������ŝ/��C�u���V"JC��z��	r�߿O���4t�P���o���Ӈ���͛7���	;v̔%ƿ[�n�Ə?v���Wq�i�id`h�o�	��
	!�D�.��0���Wl3ta�U����@�ڑ ���_d ����t�R�ѣ͞=[H>T.���>|�T��ﳳ�E(¶<!h��ի�7� mm�m[��X�`���b+/���$@�M�2EHΈ#J��ԩu��QH��_-���]~^��܎�݇]�4�ų�ReB${q,�\B�%K���o߾���*-OTp7�5��H�۷��/ )�+W���n��'�����ɳؕ*U�޾};q��a���;9���hS��h@20����hƌt��)��㏩E�%��@�AEϛ7O�cǎߜ�5s� ���|ҐU^CT��@"�U�VQ�={~:��O�<��$�6�g��1�@��������ԵkW��,--KΛ0a� �G����{���O��j�_>���J�T�IM�\����ӭ߼����|^U�� %,%��ޢa#J�W�^�ꫯҘ1c�&{k�fL�1p劕�||}*��*L�d��n�
��5����Ґ��$ =߼ys;vl�s�☏��޽�Ο?����E�gϚݟ���CW��W�|!��ѣG��G�ӦO��E'�4������Ed�8�<V�X!�d��'q ���_����w;z��K��V����/�~�:q0D��4n<mڴ�l�t^2 ɮ888ЦM����^�� i۶m��w�^:q��B��LLG&3}XR�J�mY}}㯾��'��,���B�(�������I���A�v�Z�������f�f;�|:�CFzF
��ix"!�`����M�����f҄��
)�G�#�^PmFFF4�|ڷ�������: }�4�뱄H����t�̙I�.�/%_f�S���R�q"X,�����B�8p�v���}�d�,-OT]��ݘ��~�:5ukڊ�⢨;Q�2ٍ'�ԩSG�Z|}}���@�*偈��?�����=���`[�����Qx$!R���H����.ԩ%�,$R0<~�xLj��K.��q������'z���O"�DU-^L��z�ÿ���jQ �ᨨ(Z�|���1x�`:{�,���O0�-_i9����I�G���A
6̮���#-P+�+��׬YC��Wy,Y�D,u
�={�����o~4pP��<��0=��3���2�/��0`�A����N �����`�֭�2��R#	ez������w�� ,D����RWv�����pvv����~������挋�K��J����p�גQ	�[[[���/ń����C����_����ܶ}یѣG�������B�a~����V]U�POH��d =u�T��������v��i,�� z��t�[�n�V-�����˗�����{�s�C^�ĉ�k��	#F�8]ZJ�z����~���?�[R���t����HB>����[$ 9z���Dߍ����`f�R�͇���j�JG�!M�^�x�`�7n��9�۷s+���Ρ_�t��,OOOqL&��o���6�IK*kQuHű��,�v{��O?�s�Ͻ7w�܅�V�=��y�gSϓ����[��#f���t���9�{����޸�����#�y0!,�-���w��v�yI��l�)�a3E�O5�
��\������9�����>}�t�_�rK�d0�[�lљ���.X����J"B�N�{�ZZE�jE���]��NɃ���u�x�&�A;1'�Pbǎ�����9xǮ]�օ��a.�e����]�[ᷜH�!M���446"==A���t>?����Ρ��4JKI�L�ZL��]�D�
���mۊ�F���NY�Y�"""��0)����:�����paz�d�zYO__�KOM���22ҹ��s4��utuɈ	321!K�dbnF)ؤ��$$F�҂6a���͛"�ׯ_���@Թsg�R��_g_���l��1����=����nyH��Eݺdja.^G߹Cw��!b%N��-6�}F[G�,�Z�m�damM�L����l�J�����4k�L,��y�f�1c�,���9�wÒHU�������̄UO*�
�d� �=I�ssr(2�6��Ē��� ��}C�a2�32�F�� � |i Ղ4UdT$�+�VW6�b�(��g�d�R������>w�z�*>�`�C�Rfz�4iL�Xg߽!S�F��BLR���1�����J���dmURW�l�M,,Ȅ�Ƥ��v���ԫ`�Ԋ�����[S��zt7"R��2 m�;y�$���P�F�J��M��>�@'(0��,**�	쇪,�sլ�ͭ,);+��X���>\���H���ۓ)�ĸ{JS]R�#�@@(A��������%��� �Sh`eef*���5޾Ff��
�(U�"T�2��;�����E�i���.Ā���.2�\n��
�����p@��!.&�48�q�|wYR\�6�Lҽ���j8v�!:���#ޓb(8U����E�JeV� ���o/�]T4R��z��NBCGd�9>),�~�&�w�ok�$BDa*� p!���2VV��
���z���DR���+���C*K�;H�(����]�z��=i�#�eee�rssuIE�ѫUG[tv�V�*�ŧ��r�X���e�7��B"�R����	\���i���H�$
33�KZ��
�	��5�2�J�#P�X̓u� D*���Z���0EP/v��aU���EG`*�
CE���!�^z��/u�MhWͻX$RQE)%��Ջ�)[;Hv�����ui�j{1�H�jhTAA���ji��R]�U�^k��K�e ���Xك�]�T�p!�����7j� L(���S����%tj���c0����Ҷ\�t�u��oCR ��t���rp��)8�55���XD��s�+=(����`.
˭�|�����%�zP�l/��efiAV�����>S�c	IM���lB��+$1"������(��pW�W�t2�D����RH	�u�O07
���	H;����M@
s-333���J�j�����ř�������kk���--)eg����f�i�f,��Bfmm7�F)oT��y�G�p,NH��kie%rN�7Þ9����А�7� �X������}��Dl�ƵAb�����K���qall�2�H[qGԤ
�o��Ƒ��69��_�NDdI��� i�֢�ȸ�EGS���� %O�����& �-�9���`Krk�tx@qw�R�vԨiSֳ�q�VI5�� �+��ͩq37���R)I�5N���0�H�S������A�96(�?Ɔ��mM���gR4K��m}�g213LX���EIjʔG �˖mQ}V 1!&��T�V�����ѲF~P�N�w.0�ŚS��I;"���;�#Ȝը1��+��<9Y�Ę�3RP���.F@�o�O��bˁ�a�D��.u�f�����m
2��^dgk�gÆ�a	��������`)dM���@̩�ݽ+�TH����PCP_пy�5�%B8��1D���F3q�j�?�M>n����*GY�W[����_�5J;��!�/Uٵk� �PE� +#C<�h�KI���\�9�81��_���Ey�B�T� ��@�q�xΦ�ɘ4��ҥK/���.\u:�l�"��H��)�ԩ�9�b�n�Z�6D,�-vً�qL]�� ����z��6{b�����>GG�ΨH����w�+�TU�PD��#^�)̣��2$uղe˽�7mo�~���z��AOO��7lؠ�ſ(����N���q�*��k,�^�p���k��	PE�8b_�zu�/����O���8?��#��P5Iy��עE� ���ev�BT�;F��m�{xx�D�ˇ~H{����%Dq�t mҩS���{p B *(�8Զm�&�bl(A9;,��-�P�^Q�K�9���9 �ݯ��J����!~��@A�VG�l�s�t�j����{��E��L$T݄��(��-��K<Liu�"!�Fa�X�a��� ���Q+���ǡ
����v�:y���Q�`ذa�.9(�����И��pq�U�(��T��@]�j��n�6b�-�C$�)ٷwE�D'���{ف��DG���H�F�mHLU�d<d �1�T����L���;�X����ԧ^��-�Yf�*l���+������>��3��o���Ġ����6��9s�C]�k�.��W�zC�y�2�@J�\��������]���?�]? ����w
��$�"�,����~}��߻wo���ʙ�9�M�Q��a@�Ã���@�-�CMA�e��EJ^V�����Ǚ����e�)��D�,�`����|���lе���ؒ#G���)�"�Z<��lӦ�����N�ܥ3��S��������1͞5�����°��y�Ӏr��ׯ�lP���jIy:�U�Ư��^g͚u�6�1]�HB�;��_0/w�w�^��Q[U@JӦMkIy�B��z�:�f�7�C,�x\���nL��b������q��Ӊ'�ɫ_�Ư�J���j-!�y׮]�YU�bg)OWG��Z�}��O��,/�N�N7|}}G�]�u��I�3g��}�� 60���C_�.��f�4n�����q3�&M�4���y"!"\\�������޳�)�Xǅ��K�.��*�n��`P�� �Q�yx�(q�RUUS�	:��=z�,V��q�i؍g�� +�׮[�N����?��aRǈbQ ) J���TLyR$}��Xn��j�HkT�� O#G�\��>�;M�����B�Md�2q{���ddf��+�/�i����X��Iy��HE�UR��� �>|o�~}}��3���Q�6T�ɋ����6l� f|�ƍ����	�`V�I��q�ʅ> H�6������|h�F�.�#�������~���;6n��s%PaR&�et���0��#F�x��"�Ҡa�J�_*U�It4�����.��/��6nO��e#���6c��^��H�x���D��+��t�,�y�"M�5��z9|�p��5k�����I��, �.���[�N�w>0`�pX��W�&�U�X��Q��`��ܺu�S>�b�ᙳg�ZUu���aR�վ}�_��}��Y#�$)�l��T9K\�r�Ad��077�w>4�������KG��֋Z�R���n�L�:uk�saaa���C�����\ӯX��GD��+f����?��		Q����fMY+P�:���<�s H:�:���*�(��>�~�j�ՙ�W�.������ǝ��pL�9YQX"�+��:t�@F�F��y�B1���7�/ER�VA233e�6o:8gΜV�yL����	�.]ҕ
5?/�HD }���!o޼yBxx�KPp��Np����+�z��)�\��G���bŊ�[6o��G�^AAA��U����ܛ��w��駡C�Ng����fWgm�j��F���ү)*2*���gz�͛7O:u�T?�/u`��V�U��}�1�Q�F�����������?����Y݃�Z����+R�HD���gҤI�����ݳ���_g�m0]���Х�ɑH�G�rIM�4�n۶�O}��Ycllܦu���G�����ɒ~1N�N��GEE�:}�%K��]�r�ۙ3g��]����۷���G��%�A�K1�X�����Oe��D�v�7w?4y��W_}U���)Vn*�STZ)k�R��l���ע��Rbbc�������۰��x��n�>��u�a|B��ւI�U�o�|T�_z.}o�b#,�v��mmm#����jѢš�-[�s��zHLQ��h�� M��eA��Kw F�[]��&O�G���n�~���p+����s�εd�i�4!>��<En�����Տ 	j���E#^]M]�I��[Y`���� ���D&!��u�@��c��!Ӹ�^S
�7�m���i�%A��SeP���K_4TZ��ݩ{���lv/�DGG_�����9�B���i��i�V���\.7���4B�BV+"%���������Ke���������D�Ç��{`! 11t�ʕ�;�T *S}���6�ɉ��O6l���$d��di�:�B��\����i,c��u�3�h��#ϣOU�2��GE:�qi~5��#�|T����y����&�ED-!*�ZBT���j	Q1��b�%D�PK������Q���~��"�|M�Dz�P��oL�C��[�"����~��8�"���ѝo�c#?�)��L�c)p�I    IEND�B`�PK   ��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ��X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   ���X�� �f  y�  /   images/96fabd4d-0b16-452b-94e2-688cfcbce531.png�	TSW�6~q�i�2*VA �Z*((�'A�0I�PQڊ"��"2�A@D �A���9�s����������f-���s��g�g?���^��ݕ˄�A����F�<�-Y�X�����_>~K��/u��A�����������t;�d��y�����)k�h�>s������mĀ�0m�j�;��k�w27���$[&f���tt��,�ｦ���ݒ�_n�1�`�=��k-]|�!so�O�~oy����B?I��l���K=�w4��؉#�[^����c�}}҂#n%�@�'�M}S�L�d;vg�|\������zƺ�WOڪ��g����VW	@*<�6++KK.��6��{��4紧���;�쇿V=漘5��L������9/U�c��r��;]�[�Ťk)�zj�]i�19I��DU �ƻ�{
!�w(;\Q4�_v��ͪ6��![�V���1���|�;����0�j�t߮9=X0�B.���L�0�C
�17��p�d��ۉ�� �n�=]>�����A�oVtɻ����1�Nj���v�.&F�3T�gČ�iL��S\\|����7=5��SK�����,�2���؟=���/ʖ��k�޻c�ׯX�p�@|TozƬ�N�Q�TcIx��z��j��xd5���:ﭛ�_��cz����5��V���D�Va	-$���E!����Z�����n�\6�^{�-��0~��ߺ*y�MJ��_����s�r���0�Y&Q�wNउLL��V8���@�%]�A�?���z"᫇�\|G�*�ς]��q�����"�"&"/��M>&n{T�=���j;��{#�-���~~~�ѕ��Fd�UD_��a7�rQ�2�ۇ��.M�H��-��y29�H�Wwg!�
��YW� �ѕ�=�QV$_?�l�m��7s���H/ds{W�z���]��Z�w H'z�S%\���4����_$����Lz켣���y����a����vD��WU���u���#0�O�qb�П9���!�������@!����^�}�{�1�sN<rĂbH���Y\n_��e}�NM�*l�1׀w95�����k�;ga�<T#�B_��zu��X���|MPb�[{��O�%ot������$�u�B������)ڛ:�F.P�9����3�4���s���,�D��Y�!I����I���0\��4�����2ښF0�K=83�jLӐ�OV{�;T&���{6��mr���n�9��2�fq'.�ZҜ=�l䣪��5��9/���ԙ�6���y*�w��,+%UF�lr�M2�]y��]4Y�)ˬ�ޅJά�)N9]��� SD�,���.����^��<7��]����))t7����|���e���\I⤌�p�+�4�m�!cE�Tc�ۧ��O�����`���4��BO\9
����NHk��<.Cȝ�#i*�y�YMMMK�,9H�l~}.]�c�����86VY�Q�榆�,���\�Ǉ:$bBU�Y��A�C*�dz�gHp�x��)q�8�;[� 󰱝��l�W����\l�G�.��+wI�l}��v�;��a
�Ӎ�Y�wVA�x�˾�h��&���@{@����ւ񕒜9KF
�-�:�U��]�V�ç�2�ko�sn��z�ah��d)����
��mN��e'*�[�rFXOX6�[�D�ħ�!L�iG����I�P�qT�G�}}���{o0�N��s�x"����Y�f���]�<�RdX��~��cz�Q�t9�H-tRv�H�N��=cn�a�f��fk���[��?��B�eΉ N�]{��&D������!]��Z�=q��o��e�~�8'Os�{'������r2�p;�CD�zݽ'i������܁�---�=���>�|� �"��5�͎�7B�=[��_�K��΋7�d������f=N��s�����0-]K�S\sXˁP\uz�����UЉ���4Y���xM=�yp�A�s	-b��wn�ϻ^n�34W�pc��Y2rEA�.��`�{C^���;UaG6hsl��)h�(�Є��G7U���d]266樫m��ކ������=6z������-�Xw�a�z�Rt7� �$�](�B���-��s�G8��YhU�� p��r��v!(e21���R0��~��z��F���VnYM����љ9�tM6{�9��iͿ��*�&#A�o�g}�Ɲ�q#6VL�┘ds_��$J`����y:o `��/wti1c��?r��m'^$m #����K Q;����ֱ{��1;J�uC0�0�{��v��h'a��a̧QJSp��W���=���{ ������q��"-�l6ȗ�2  H��f9V���
�K�ȋ@�h�
 �d�W.��5r3�{k�Ó�p'u_�"\��F�V��F�nz���CF�����}zvNMu��x4��<�5b����Ҩ�,ض,���R��˗/�2^��o�a)�\�X烠,��O�\	�����*�W��KJ���a'��d����H�4�%�U�Y_��DgK�TlB�m��E���iÅ]�Hٶ�h]�� �T/^$R� �d����X��\����^9ɪu�uM9�![%� a���M0fJ�3�:a�f��A�8,d��h&���X���dե�fҔ#ybvz V)��R!;����2G��[�'0B#Y4͛s��ϺC��@��l����N�.���� A�b��(��g�H����\U�r��ٺhONl�Y����K:�
��g��ӱ��X��G�Qn�Q���Vu�ƾ��0�CzL$�%�j�M��tG:��|�2g��_�����~z����' ���p�R��X%V7D|f��fx@^�
Ev�9�jN1���v�Td紊(pO�#���sl�T��c5��B���Uy(��&�)S��&�\�$Mw�s�zn>�	ZjêkG)��=]��wX��JQǖ��������nE�?@j�����}sa�
?ᘗ�i"H��	T7o��+�6����(g�׶s%[����圀����DS��Z��\���y(Nz�DO1hXaD�J8�\�����;w��������,É��6W�i�����e���|�>�@�	��6��M���WC9ɵ�o�3L�@a,,͠D}*I}��4c�r7Ǖ��cNZAn�Ct�ׯ��}��u��9i��
�R�B���qW����Y|��i�κ"��ۦ �]p�o��	HJ�;=ҳ��8��1�*Q�t������p��q�^9ȕ�6]����Ɯֺ�'�1tqV���"(}��H��l�0��h�0�5.�RO�_#�#��gPrgpH�f�z��`��زT�c�T��$1.��Y�( �(�t+AzvI���)?�hD|I��Q( �
++��9G��G�g[F+~����&�К��f��1���g0���G�D�t�jDG�����E0��p�S�}�]��-oQ��=BPbӥ$]�n����E�x�E�.�R?�Y�CN��k��l	
X�É" �XM6�����q&;�Z�`�������D�~w	4��<q���J�����uϩ2!���E�5��(�8vu_�q�qL��5���V-; �+
��cb��03�E��w@ˇ���1�̠�&5og�;8��9��=�N�Q��(�q������H��9 �)��|����ŵ�#r��Ǉ�z���s;�EͿ��-�PN[���Q�۶�:xF9Ҁ�
��D�x<ݲlf�9�W ��xމ��=)�<ǀU�_p"��0T8foZ����Ć8�' �U����3�ј]s" /|ŵ���6��i��F�Y�h�֊���n7a9������l����52�X����zw�0�T� ��ӳ���K`���/9����
�N����
/ւ]q~�4�ڠ���I��R�zU�R�%>�`K�e��@%UI����_������FI#��o[�z#9oҽ��w4h5�o,$�K��úW3=^0��b��'��պ9��՛���'��A��[8�����֒P���\��
q:*��WO�����5�Hl+К���<u��l@vyV��B�(��A)�ưi6���WC�����6)^�� <�]�T��:�E�y�K��DϬ�ǽ��5��;��_�ѳ��)�N�Ɗ�`�p�Ig�(y�n ����|+v�S��J U��)�q���g�H��} `��\n��;�C�<�����Xxt���,1��;eJ,��-����ӢI���^�%ڍ�j�oŵ0�mn�$�ܩ��(����wS��QʨfĘ%uf�t�a�ujR2�H�tz�W9*3XSQZ9�7A��W�1!�?#����Z=� T��'_���vd6��`����Y1��y'��;�'C����r�[΂̉FrD�:�(дTm�ZUcBgᓽtV��%�Ŗ���m�����55����mQ2�����sYuM���~B+�u?���=��}"xl�7i�#������I<=��.)�{�z'�[Us@��a�q�Ғ��Y[Q����I3Rr��D�O�ƺ�61�LZ�<|E�Z�C���2������<F�`���F��֚��N5خ&�^�w�	U���:��٠�Żkw�ZE�\�ʐ��w�����)}�	�j)��Vs�ۊ��X�ЗFRfӱ�3-���{�zb���Zw��=���͠���(:�w��v��qqX�M��|���-;������K��֖K��I��YV� Zi�q����c�|0q�l������Uº����4@�5D8�i�����6纜�B����pŮ�D�שr����錩�<�B�Qf1t���Hm�޴j�e� XUL�b�'\X}��O�
L����i��olA��(�2�~$Bc)�-�9#P�����{3��r�t��mS�#������Ps���D�΂��h6���ޓ��y��Zzv/�(��^Lb�^����0؝F�Q5�3�r�ӏY�)��S_���ꝰ�m�sCcb>`:^�Lc�b�7:ekK���=Un#/�
�zk<\Yv(F����X!�{J�����zW ��t�s����\ˎPF�/�&�(�&Oh�w��a�<��6��B�1/�'��ş	�~�rl]���0�����oA/i8��lz�E%na^T���dd
Ut^q(���M�����-�̸Q:bA	z�[C���;D��89�0�zq�!�4g��gf|uw�4�4$��.�I 4�?;[�Y��[8���9S�'�BHjH����b�pؚ�����T��1.�`5f���KI�YWԹ}�2{�~b#A�h����2�\<� �20�VۖA"v�?7�ۃ4�"��������iP�p�"@�a$;�����}�*n��� ���d��-��'���|�漾����u��ɬVKJ*�I"ܾ�Jr= �v!n�r�!�Zܸ�Q���D��3+'KnII�����(Зc'��1�"����e�
�o��0�p������d�.�)� m͟��H��#�K�9�%��zO�nS���Ld=2�1�?���<k� \�������y�����%����p��� �U��[%��g�V,�¢��m�Ŏ�Vg�E�:f�W�<ȭ,"Qs����ÑFk�څRh����9h\�*3����������p��t��|�ۛNZ�.S~;+��p���bkc*��|F!�=*O�M��nM_�B�����󲹎���[W���tC�t5@���d ��P0������
*<�L�;U��M5���q`}�/C�p[�ji��kd؛yy�C���`��$�S�[25����	��c�Q>�h���\��	�t�	j�{�Y�5]�<�y����5����� l.P���,�䠔�f������+�\8-�p�-�e?A�b��d�"�(ǫ��{u��#�J6]���pݵ�}Z�� չ.��8<�b[�,�&�K�`G�+i�ۍU۱��&�'�-lϗr8iP>�A���P軜"��Cl�-�ध))��+�A�͢�;����,��tfm!��Ť.@ڲA���y��w	p?|&��PG�&���ښ��)5�Pɴ0��&��r��}λ e6)5f ѪYط�� �0Z����p{}��v��!���[гVШ�y!�;hY���lȲ1���y���������"e~����Bз�M��:K��������էxJ�3�Y��G�WB�@��P�IF��L83�cq
�֜�.*&����0�lH��Y/l� m!hi~mry�nZ�����iƞ�2s�{�[8#]����&��2{C��y
j���h9
�I��!�f�6�O��	�=��(T��^7Y�X��i�sQ		�:��AW�ú��d��t�v�%姶9�B��ŗ�}����4�~��s�) �K�,B�_�U�?������qnv�m`��ڠ⎱c:�+�u�&���&^k�MP�z S1�w��jȇT'�A��m���|vw�jD7�@O'n��o�VE&�8Fy�+k>{�84�Z��~����������?9�l���;��^�����џ�X��	?�M�!Yǿi�㭗�s���2���Xq�R���Z�^u� �hB�}z~)��14~��F(b3�\�e�M��W�p~z-`|�&��َ%�X8W�a���9�'@�?m��9���Ț��{H�A �-���7�PkVw+ڤ�O���oHӒe=��v�%�5|F�CŬ�ڒ���-Z�l���=�A,���ه`��S�X��<�ۛm:���G��}�ټ��=]8� ��N�e`IU�l.��c�hp�{����e�d�Ѽ�A)p��[rΕ_X��W!�����W���V�
o�ɖW'r�n�r22�Z_�o����<ӣ�ـ㇭�(ہ�ey��.�>aN�J����3S36t������cT�8�d��j����$P/1�P�Sߩ�4-v�'sȮ�CB�PMj?(�0'�����*e�R�a�l�O��=�l=���I���
FYb�)K�sO��t��؜�/?���d��G�il��ϒ���䲟Ӓ9�2u����,�E��s���6\ÏR�9���}S�{/��w	(���cЎbG,��/猋��s9�+9��W�c|�{�B�D�N)��>@���:9�T���s���J�ka= G�P,(�8�����^��~�I��f��ps{��w�����RR���0&y77�n��亨D�iE��7�C�i���&��@u �:%I�� 2>ݸ-=-w>���I�0ψ$�^����LX��x�3��M��(I���@+�J�>����Է
�Y�}��wKj�9���z�Ϧ��x�շ�2�Bt���
}�����ث+
j6�6��!�#�c7��ى�YΏ=��څM��*�s�������[R��쎇�:�Ŏ8'���|O�w��ʋ?���z�H�<9�:r�1*��ͫ�Z���K��&�{���~���bK���Ǣ���o���t��}��I���~���r1��M��BC� ]����z�s���4�� ��z蜝��J�L�}H�5I\p�N]e�U4CZ�f1��cvGv�4��c��B]�i���p�->o.��fWT7Թ]�vmfˏp��.�����I��qHPCj����HS�'�zqv�.ǷAj�}aF���J��DχzAW���n��j��9���d/����;3�j�H����<QA@��m^�΍�M�H3`�}��I��̦��ר@�J���ũ'XW��Y{��f�|`�=ˠ��t���-�2�r�`�0���F0ڌTz�Qs&�9����T*���A�i���=�$��P�ej�������|dl��qkAzzd�>�tU�4(Mk�48I�4o�Y��y/�GWg�]�Vp�I���P�c��%_��Ž���&���$��N:�ň��T�f��x0.�b�َ�m�Bo?||�l��Lv�fsj���q&j�2gaFeNP.�3-=E�PSS[Lu��el�x�U�G��}������e �؃�<w�r{g�-�op�q�����p��н�|R�*k��܉�Re}�n~�.](�b���"�7��΋���?��.�A�n�ºu��Gkf��0�ys$�ʻqL�UEa:��^_,(b���`D�ǰ�@^�M��\6�V4�xyqJ�!��Wp�R9i#����%��Ka���?�q�{��� ��魷�4�[����LQr5rb!�gÀ�n��n7���RDӅ=�,*㤪Ho3�7wgL�|.�(�0���!7U��`@|�e/[@'bz3/��2�Ҧ��ϑ��Nn��������j�R�c��p��>q��#c�hE�=��_�@�Ϊ�Jbe�?YPn�R���K��Ka�$W���­�I@90=pYP�+z���ƹ$Q�����J̪�Y�Kf��Fֲ^�dj[J�fC�K�+-�����:r�=P�r����Ĭ�E�=A[�eZ�P����]��4�pJWH���4LS9�49���5)5W>E#~W�A�M��ܡN�׻7UMM&�>�P-��X�0�q*��~��k�'��)��^Ajj~�D����TMu)Y04��4�`�aq����Lſ�D���R*���rnQ��	z&P,�=�������{�#���H�$b�@���&gS������1S-gf�Dʞ�	���]����	�������=�d���\�?�n�����������������������������}�.&F�?i��]��@��=�ֽ�Q���u�e�˙а�K�S�={����L�ym<�8�+!��B�qO:�;)����C�#�7j4G�$�I}f�M�K���`eb�Z,�G����#G2���F�&��뭣�X���!q�挽�~(��F˭�	�k�*�����Oss����N��9�6�����V�xa痼�����h%��Ω�FM�P���ƐK�ǐ����hh��Y�Sk��Sr{�ݛ{wwe~�c܏�n��d|P�b�Ӓv��2g�<��}�NIL���=PlK:�tAe�@��"
�>�u��3,�,�9)�QnsN)"rʧ������gML���ه�:��z��?��r�������q�/�i΁�w������[��ឍ�>���q��7�{�_ޘǬϊnR	PX��P�;��ҕ�5��+*�eC�N��]��Uי�{Ϸ�^�s6�]��M��-R&�:�7��5%;�F��q�2�e����%>����}��,�#Ci�}���K�����K��@C�i-�)�c�=�T�;��DȐ�9�aR���G�a��C!�M�N��f]�+�\�Dy�vf�BH��$�B���ֶ?�2�);]Nz�KIj��A�N�ZagF�r�B�i>4��?zo��Ջɋ��v'�F������
�Yu�+�ϔ۴�T�MLu��qvf���ʨؤ���x�>�Ŭ��
���{&�Ns�������� yG�@�|\\�����sg	��mf�ŏ��Ë����@Hq�G(��άoqs�e���h2G1����K��GK�Zf:�h�9��b�r_�ϫ����l�a1��!�8�}gggBL��p]�&��o����dd��O��o!�����	����@>6��M9�l+�R�r���t�����5�gI�Jc��������[S�\���X�i��
�M���*؜����
ͬ����
��DV�2��Z���di�(Qa��|��+�_�ϑ���b����:���w�����
c]����'��`��8-D+1���D�l�Gu���t������Kjy�ZӃ�}G{jz�C��`{Q`��%��x�.o�l� DX�r���	�%kwӠ����?���͇�z(��N�2�A���j��~�]�r�o��SU(/�'̤�ncA��:�O�Մ��?�*[_����G�we������o�v�X'�
�p�W�d��[\ބ
�( m���:��g�c
y�Ajq���%��M<��'�D����@PzJsV�:�^M5َ󯣃U	"ZZ��*h#��"���V����+)Dg�!��h3�	|˸����0V�2����*~����KJ
���R�k�7݅w/&��W���!������);!����
�z�_�m6�H�Z_+��n���λ>"c�|�.T��~.�kV�
���Sn�ŤƗ1�m+�Gsn/_d-7�R~9�O���m6����� B[�W]��-P�a�"�ٯ�η�a9y�u��-��6�\
Av���< ڴ�)WZ[F�y��4�T�o��b�_���	��#���ԻF��I���_�M�v3�k+ hծ�ry�ҽ[ѓ������n"Q5����ȷ���`�5�Q5���*��� [1�?j߻�Y��'���%���m!�91)	9����k+�P�"\�[!�{Q�������󡽚��MX�5��4��y2�G�������شC4E%��'�W��dM��J�Mc����׈ VΡP�W� �y�J�G�,fm���W��M����u������9���+���NP~�
A�G�w�$B$���)�������\�OW,�p~�8_⓯��_������_S�(T*�� (�%o!W� #.�R���s���t� �����s�x_����A�'`!���L�U0f]��`���J����H+㚗��w���S��.�<m��$�L@��J�t���L�"3��Oa����(*�Ȋ�����&����Z~��p	Xi��1 ��o�C�_q&���tij"h*[P}��FezO����X��r�K�׾_|�ja]���ѻq�YOц���.�:�A2N%�hVs��}�]����C��T:�˯*��O�7\�3E �(�ׯ����c�������t@�D<�^J'�9�Ci �<���V�G���ݹ7��U��X�������j@y���`<�!\��^� �C��'�'L���,�OM޺f�B~Ś��?~h�s�\{��|1��,�������pqۨ�H��0N�/@�t��H
=v��������d�"���[�������߉�K�|ʎ�?��Ż�F �EF��o��q��0���x�����5H�2�}n��Qa{/��R2�Ex3�>�+76�{��͡FC��ٜ�����2�U�?�/�����Ĭ��aS	��mF�N@�vgtEL���7��B��������� �]����߽�;����Y_��qtnػ���@�j6,�&�cU�ߋ�'^�k7�s�u_OO?�s�����Z�C!Z�Q(/n?���ۡF�w�&�nE͗M��F �J�Hg�{��G�@{� �ٺ�3��2�c�V����$�T���~c��@���>�6%%�0^W�r��k����ZS��8�oK"��NI0�`�ay�g��Ъ��o�}�n�\�6~Ϸ�M�!����Um΋i�3�+K�c���ʓ���������T��K
�廇\Y�;�����3��-��X��쒁��ݠ��������� K��ļF��l�H[�vgj���;-�(�Z��˩��wF��b�O��t�(\�14~9�z0񋔆�`���hW#�LQD�y�����N��
���o��maN�,5������6�@Z��ֶ������F>r�?;v�I�՚��|�#̛�M��J�
yvƆ� Z����L�]�l��i� �{��z�v�����V�N�U`@j�������s�d���J`���L�[Q�\��Z����3�B���嵴�g_\Ӻ��������hÞ�وЪ�H��+Y�<ˣ����$A��{�ױ��ة4l ���Q~��I0)z��#˿V��n!�����d̚���4�G�k�>��Ą�ؼCQ<8ǅ�����k��	�P�v�p���FLL<mwww���
�L!VXQF��-���1���L�]�r�H��5�3-h����0�.�5Qr��~D��Ԯ���դ��2<~8'9�����d���qu�� f�y��WA"fH*����w�&��.����s��!���ҒJh���ҝ/Ȼ���nnktuu�g^�#��_/**:ii�y�E$�Uxb�S�V�M����
�� edd0��>uq^���`�S���0�1!1������G�L�ə=[5��笉�/�_�bl+�<�=ݥa��h�F쐕��W9�p`pql��
㔞]݅T��6A���cD�HL�e��f@Qnb/�콙���i�)�!�(+RE%����^���%��4Co��j�cZ�OƓ �͒ͯY6W5�V�vy�G�?�Lu"�֎�y*��-4ճ�32���W����H����Ļ��&�����Ӵ4���w�?o�`PA��;:ć9(�#{wz?f��h~���
#�j�/��a������mll��!�~��.c��[RɕA�Lv��v_]���jޔ�������y�ӓ�!#<<���f�u�N��ț&Ԛ�e�g�P����X�)��4�_�!a�F���>�J`NS]���79*'Zd�	����Y���b4Pv>����������Π��(88�د]Y����v�l���.��LF~�g�_�g"��]L\�Um�	��������L��7=�Z[]]���zݲl/ě"I�I:4����W�^��[=��X���'E�b��3�+ ��V�T�j�_���N?)���c}���p��H)"��x�ԩ��1�'���J����Qߏ�۠P��
��l��ɧ����Jt�2rժU�Zr%V��°�����'m e�>�s���:�C�{��wQ���]N��	i��W�H�x_JE{J�f v����������>��Y�)fć<a��(�3�n� i��6�b0���-*_Z�����L��kaD��lR6DP?<B��mI��5C���xQ#=���. RGc07I#���*��̞���-�Q���>��(
u�А���^&&5����3^���Ky4@����D���c��@���=k�/_�4=��[v�����Q���Rw�Naˁ�,Đ�^wf����&S�<�.^L&���i�ɼ�� 0�$Z_e��]���]tfp��;�HT���5�t�>�[���Ei��#��.���(/+��~� �w>�Ԗ��Hۜ9�@R�]:^� {�d	X��4�1И�B�5��I'�������X{G��\��Gܲ��+
[e)})J�|~t�p�ATDdd�|�,m1L̕�N�j����d�j9,C
3��[�̙b�SB����]/^�8mo��^��99]�(�F92�%8 ��T���]�� ����ʾ��m�+<��`�U���3S�/F7 ���?`hU ��ddWWW(S��C�2�6e���dV���T ���Yb(TQ�=�Au7����툧�e�ff��U�ώD7�{�	����j�5xO����pU���(��熝�K h�v>�lc3u��G��`2ГYY�1�K�SBR�P���xt_Qs����P���� 1�Ԏi�=B+����x'���
��#�1�]u9��b�mB�s�$m���@m��'OΧ5Tv����NH茏�$�s��Q<}�Jk Fh����L�u�2��1\MD?'���m>$�2P��<sr'yy��϶Q��4�@S` �*�"�s���'��3�)�M���Qvt���r3��K�ݵ~�I���m�,��cH���㴭����{�D"�B5�l��)2qqq���7 ��D�@|R�V�]�l>;ҥ��W�*4B������J�B��R�v1I �j�ʌ0����H��%˭ꦬ&GE�$�#����c0+�<��%+}�w}��{|e���T#�Eu���������⎺����I	X�?
�	�����5]�'��0��y889��O�i*( ��Ў�	�5�kIꝌ�+C:�Lʹ�z�e�ڟ��@@� �XP\��)�A���T���Mh��l�� e P<����#0�?m)�(,Wn��0s"��̍<���l9�BT���p;��A�&SR�y�f2����������u���!��S�"�\"Q<3��,���A'��:б�o����M�(7ZМ�6�цdp�L@��Nar�9���BR�I$��xG��1��,��i�^7 vy@:R8h�7s �:Wr����cE��y�e�>q�y��S.��5�;/+ �OĹ���j���a�n;�]�����qfgh�v�� @�%d�Aѹ	���$��E�]<I�����'oe&2�^�d�=I��T��x�g���Hs�pQ�该21��xV�i6f�E�����ˍD��"a=���Ǡ-�*uo��BG�,1�_PP���~󚠄N���!"B�Fjr��N�|���Pt0p7�u+�$E^Aa5`)�]P;�aeb�RS���u^�}Ro&�i���EBi����s�+8X��+B�l9��:�:�'OI$����J%8SZ&	E5۹�?ाLBL(�e��i8��#c� 0|�4�[��� ��
����n[�-�ߣ�0�@��Q���R�*�ng2�i ��=�|�_ ����1A_Q�O�'�,-M0\�������ݻA�Y����M��D����쎕���&��清���/��F+���L��N�N�Nk�,--����G}í��O�4�=P��~�W����b����ک��z������9�&}}�����ޢ��;���;F��23�{�XR�fW�ׄf$xN�:��ȶ�ZO�	�#\��5�5�Zx�$�F��Z�Ύ&E�\8��/�ٔD ��ڀP֍��XP�����^��B�-�>u����A:��ҁe��I����EnG�b7���HH����h���G���roNLL|���r�`������_��i�SQ��K��u�{�,�<�LN��&��&��=�O�@��>^��3~Ƞ����quD�z���ji���O�y~�hr���;��&Xao�篵��C:*�u�}��$a��<���/_���y!�6QX����ud�&m��REEE���M����?7M }w0O8��,���mx�>d��a��W��;
��O����jۣ�XC������8��sF�u���Z\'��E�4қm�9IF�Տ�@3I�o�G�����#-3^y�GQew�p,?�$)�\�?�R��f.��F��J�:L� �_d�7\�ag��|��u�C��l �<�a��k���ƺ������5�6�ު�ݱ'J�.���U���?�AxC� t��m?mrǋ�u����(˓�^gl5UIA�mf���	�?b�)��`g&{��t,����1*�
ᎎ�! 2��I�Ɩ��&�l�̤�V�v�!b��l1�+K�2�<����6�0ةP�8��l>6��>4$/.!��h���r���9�"ch��a>L�`X�񾊢t�gq���4�l�ι��Nͅ�	�YK��h�V,oHC�pe1�v�C�ձ�m��A�w�����o�\��ݛ%<Q���5Ђ��/��-E�K�x����CԧMJ� ݵ�ӫ5w�W��,:��>o]xw_��"���މY�V�s�BS6�$oe�w����{=�'�n^z���\`��T��O������K\a>$���K����S�6�*�yVI�w�����z;�	��[���I��_�w�o��_�^���;+.��m��χ��R{��@�%��!���=<��7�@�%��&�D�'�Hֶ�6�F�M^��u����:��c��&�/?�ٶ�f�N��p(؆����<�p��M?��]]j��}Pr��dYQ�|]�L��3|9r9��>p�0�A��7X�]���o�y���V�q�+%��ٽPr,��!m��v-�;�+[y��~��}}�K�1���hyz��H�8^[#dd������@�ٻS��9�`��;��Xx��K�hn#��_�� �;��ut����g@���ŗ/�o����n���o������?yA�)�
`%<�j5kk^�١9㣹�-�ʧ�o�����@�������y��e:_�(S���H�O6>�9���Q�{�o
�l|Qt�n`�����0����7��pk��n߫5
��}�a���l J�������,d�8H�����AQ�V6Bz�������p�͍�]B
��y�������̳�� �̹G��_��S���>�_� �D�η����T����I\�u��
�S<^9���|�`:ߏ���D<�}{��.��W�����t���n�Z��l����*`xy���!6�_�:����.GȼxiΦX�6P�&D��� �� �V>쇜ݬ�y���0ʻ�kUa�p� �R��v�ڐ׺�K���E�������${������zo��m�|N^����9�	�9%�����d����ޡ8b�f(�[��{>�<���90������r��i%������_�q"��}1Du���'�]yf�[�K ��;ͣ���8�2�]f����jcF�c>���������m���"����W�8�Ւy�ڈ8�=�5� ��Ȃ�)J���_L��y�N�l�S�۵�l�w��+��ϠA��Cbu�^&@�':���qq>�G��?jȤ�W,){]6�4��Y� *��V��&N����J�q��:=��?���'�x[DӏM�z��������Sޔ�{H]}j��"��_�DxG�O��7W}���I�Mkxt��Z���ew7�a��eu�M�dRݟ[k���H�o��}V>e֡��#��>6�>���ҩ�oӾ�<=�b�J$�M�K�\�Z���?�-z�]a��I�(�y37��{ץT�d�����W�/y3�
s%N�4b����t��<t�|�v]
�����F���TxA*������'X�=x�ܛ,�k�ª�yi+��$����a�û@1_AVm�~ H`�O��N�C]����G@���+@��%ށ�>AX���ޯ��OQ 9�Lɲr0�ｚM�_j\>S�k��9�|�h�I�d�����C.Z��2����]�{���E;��}�e\��L��x�!�BGy�h��s�T�'/7C*�G��Nyx��ٞ5 !�/��|Z�Ma�B����ޏ|�anT�2k��	`��_kƹOk6���n��G�V�/��7��b�~Ee�E����BC�WD�����^�ֲ�����6��{���5�������ξ��(��ln��	�D�1�)t�Kl;i�� �n���#`�Y�dz��?g�����
�
c�ྔ�/�0��/;�?�$��l	۟������ѱ��F��:�WF��6O='�k
l7��>�d h�ꗐڕ}��_l��f�����>���F�<�����u���S)�ˤ�ӝ��!��Dj
PsC醹��x��E���A�;�8�v�%�JA�d��R��
�9zy��ҳ�]���s6�������r�B�~�<�q�~����O�QV��7��9��&@���%g*����kW��]���4.��a�`N|�;�H����~��$���?�R��ħܠ��k���̗��ؿ�� �`!�,���aF.�ka@�#������O�#> f��Z�|E)�t0�%��o��k5�8��y|(�{�<��I@�w
�-X�wun�������X�c3�e�[�~��蚮��� �u�����`�ξI�d6�?)楝����@kp�Rz��Z9��a���p�n=���u�m�I�<��|J�<�fėg_��{��F���&h�=�hp�L�.�6i1�d�%$�X��_8���k^,��ټ��4wp��#�D�R�~#ZkK_Sӯ�T�!jx�@��x���N�n�j���7���OF%Y��ɛ}�����n��Y�I�z��/;tm~����ͳ��̻��:=�҅�j�oI�� J�L;$7Bc�$�"9� ����ePF���������/�i/K��x��}��ॷ��yn�,t�H�BEb��%^d�m+Ux�6�$��>Il�>㳑�`d�ʁ���Ep˩���v������`Lm�Mf�P��p�|_�/ ���\ܓ��a��jcjƼ�!tK:�,vh^Ŷ�f��E��렬-<�yp⣐m��˙�C�3ߟ��yK��лe��������c��릿Y�=@)�;����E��N��'��^��h�)�g�~#�Ʉ�yG����u�0�^i�؃���ޟ��y�zA�YS�����S!�ao�M��"g�`���P��= ��2?��o�f�f'[�m_!/a�T!>�@�Ύ�y���d�O!���yq��Tw;�W�Z�my���������%�E�ƍ��;V���^�I[^_�{��7�"�4?��K���͇5��W1.]�[�x����0�##F� <{������i[>�v2��G�8�jp%����+��L����?� ��\�>���W%owT�j���/���[x@��h��(�X��J���|^�_�P��%g���(���3��?����"��`^��~��:�� x��ڌ�}�}��ʁ�+x���A����ὭÈD��b�4�[�<��e_l��ح��^u�oc�a,�3�u�N����	�$~�XO����!/ю!��
��x_,P��.����Vrb]+&u��)�Iv�/�\���E����rd�A�L����ѕo�w}�3=Q�44���dU��F�
�8/b-��$�<��p��[�����d�=������9��^�� �n�)�R��(�Aޤ)A.o�8`v��|q�fq��{[�D���$F������Xc��O���e��߁�F-(�G}-(��	�-���hM�{]�����Q���F��4@G)�2��*?�(,��ur��Ҁq��h^�&����+~wk48uރB��{�|x5
�0�6D�݀<�Z���){�oY��DW4����6p�{z�^�y"������*EVkw��/Qhƥ9\H���xx5ۅz�.���3L��r�ǝ���1
��n	����:�n�Z])��������<��X��Xq���!͉I/����R]�mGA۠�1�j�^�	#=e��Ս���>�I��8e鰵�b����L�2���<����R��dHJ�.�^�Kʐ�/D�e��8V��x�8�j<��{q�����<�/�E��T��I}�A?���YE}���G&�ߴ".�DW1��4+�dm�>��+��ÚJ�}csm�ሂ2�� ����r���$�"�� (�
���Ƞ�AeN2�`��9B�H		����>�{�}�{�����^��?ػ���Uk�֯*U��!�K�|�>���u�O|����^������Z��OE�8&-q�g����`�$/��UJj�L��I��X���/r��
�3�Cف�[ �6�m�F�.J�(P*�;�Y��h�R5�W�\">p"���-�0MEɜ"������K��݊����R�1����&��S[s�#w�GB��w�z��p�߶�ZYZ(y��q�q�8�eu��9Y`1�w����p2Q��`C#""���1����o�#>ǳ�D��Rֳ�9l���r;�*P9� q:4�i˥L������5%��@![�}9�&����Xÿ���}Lx����<Hv�)_N���6N�7�(��^ڑM�.ܵ��뉫dĤ��ޏ���q�<9���=��)��Q��&��K*�|#�i�S�c����%����_�R��9�k��M���Y���礪�+L�� D��7��+ֱx�s���%�������	�m	7Ʈ�~@^����D�$!����0��7%�3*"܌�����Y� .�a����~E�M��`^L�G7�� ���)ϛ&(��t��|{�1�#[�,�6��4e�����z*���lI�����V֚�=��V��
�Z���K@E�u	X@�oR�&[Q7�(�V���+u�P�5�<]�����J��=�Z}턆5d������9r6����b{t�AM_;�߿��i��V�Ujxyɸ�S������ֻ������w����>�I�AG�����;l���$��`�)0b�ʘ��ϗ�T�M��2T���@��W�p���D�]T'�'�T�}����M]V�|�*L�^oj��$�Q��=��7�U�1�r�=���!�����ʈ�2��[����I�'Na���-��Ũ���٤xg�z�����g��U�7o>��Rf��j�Eǃֶ�k�y�'E���`���/_'R$��f�A8(XhX�L��Vg[� ]��%/�Lꥬ̮�T��7x禍�i�/��b��~U}���0p�&'~����q�Ĥ$�TI����@�c �c���P�_*��3���B��*vtx��X�WK����b��a�j]z�������vk�u�2��yy�k�I[ 9ΧW0�`1G{=巽�o�K�.��Z-j��U��`*�`�*ʠ�ƛ�yܰ:i %����L���]:�%�ɐ��J?
S�E	��f����,�l��M�'��7e�Ol���>m���)l������N�eׯ�N��W�Lкk�ޜ�?}�����4��Ջ����tf��!5~Csssg�����2����@p��7o�H�D*�n����B����|�1��=�o5�I�M����%���QdT�ߺ�`$��볘��$)�> �׺�q�+K֋�L���*L�ș�Q���,�[a�p?zt�Mxa�J_���6�`��m:�P���"�A���Q���{�/��L�J~�?pa��5�s?�A-���G�'MB�`��(�r���`=�C�%�I��~�q}���I��58�����In���
��I�=��c�2�;66V;C:�箏~�FV	��E��*/\�/�h�(!����	��N���( ��R�^h8m�V�Zu5ֻ���?����=Xuwa��z}o���q����ʻ3�X	�FN6�N�q�n��(����3��*��'G))'??M��7ٞ�:b�J��������\�n�u��Q�Ԕ$K����+�-/�RR����sM�� t)m�`շ�r��įC;�S����K�%�g�'=�OYs*P�U�o�Ye�n�cw��s*	@kq������G
��V�I�A�k�wDM��%��0�B�ׄu۶��:���!�#:��J�_���>Nqʦ�I\�'>H^���#�7&���t{�>����c,���MMMSA����=����f��x�Q�%����P�Z��2B%��e����6#�l�hnz�p]:p�����s�-^'�%�g̸|e�v�R&�`�t����z�� 6 �o>�Z�����ܻ _I]�5�z~q	>�C"߮l(}F��v��{%�M>Y���= �W^�t~r )^%7�֑/	�}����m��b08{�=��>������Ѫ)�:8���*�D��Dݵ:	��'���_�I�|q�̊i��q�1��$Z���� %�D���5���lRMpP�	Z�_�	
{�}gǴD4�l1�=�3�(U`��OB����S�,e�4�T��	�jev�y�����O~|���(��c�5��.�S���#p2<�s1�[�!ǎ���D�� ��~�[�!sC?K���Џ1��Y����2�E1�PU�����`" -#�]?���a��G�ېW�� E���7�_����L�� )FE�m���V�޸�)��X�:EC,�߃-���ץA'���8�4F2*Q(˴|�?��#�M4�x��|Q&zௌ�P�N�Q��~����ba--n�ys'��*}	�|��ězg����vY	�(�@'�1���eC�����8/�j .�q9�������ݤ�AIh�(��(WG0杳�Z�A�g/����.�d	�$��1�.��ԡz��@�s2�`ʳ/*�5���V;fQ~�:Z�"��{����kP�� V�ea��a�ꞿ�̿����~����Q#ӡ��򺓐b)p`�`�P�fЂl8�ֱCPV9G(���hM�eX�[@T�G8ȫB/�A�Yd���}������o4fL���4&Y�f47x�ɑb���H��A|��(˳�f���{����luEb��(�b��*�ΏP��
��=CN,����+���b��RF�+ �d�I�i�r��q1�x�4gQog���{��S�l�'�;��8<,&.}��4P&�S�.w������I�X'��ʼt�-?
Y�ܯa�?���^.b�F`b�;qaf �o=
)�x�a	j�`��� ���5�����_�	�3���u�2��SR���L������/KY�����ԪP�\�P\D[�@�{���;?�׈l��������W �zc� �جm��2�kGA�g�wy~tkG�ڭ�G�[�Y���.q�r��zv�a�:��-�:J^����On��{��n��8u�Q�a�����L�����%��V5��ѡ��/v�Y^��"hSa�Y�#�x�e�g��D.K��/�����	��Ē(Ŭ��&�Θp�s�/JpM���Ж�^�ho���R�sGǑ'�!�A�����#�=J�����c�OR}e����+��ݹ��F#Z��%g�����wkoƄ7ekdtU��q�2�*����9qC���N�M��@0u����ʯs����JY���=�B}[w���??w$ԧ?�S�iA���y;�0�����bL}�>��+K�>󄹹��%��O��<0�Z��)��~�#���dۚ��V`��R{�����jT�za>��n���l�n�-��Ź��=t��[ny���|j!�?\g�v9u���ߤ�z��V�\h��%�ۻ�љ����i_)n���^��]˧��۝���l7 ��}"_��t��7�]����mK�8P��60'S �eೲ<و�#��(!��3��u]�Yn�l�v;��U�S�"q�N�[���NKd�(P:ҥ�����n�{�\���>B�����۟5�Bޤ�+��E!������'[����y�e�O͕�,M�;Yj�GFa�vlp�U\t�(S_0�r�.r�b/\_�\i5�ф�§ϫ�''a�~x�;�E�͠���龧gTc��t����с�n��B��2���oܫy&m���#���4����z�y�W�����s�����x�@���<x��R��y��CJ�	��s^�h,��P�%���sQ[���&��G�ܡL�*tV��ǫ���ݚ�:d`�~���ߒ��d�6l�Y��L%<��������v>^��������|�~�ͱ	xw_�����D�IYz0����X�=ٷgg+)�{M�P�)�qL��A{���Dn�*���=/�caFH��J��~Xٴ�����ħ#�"~ﮪƾ�%%j��[�@'`�^����D2^��d[c��@Ѽf�e��SS�������`�n)�:&�[͹������XI��҃���vS�^�g�� BH�����j]�Ε�N�N�c~t��^E�R(O]�^�΋��G���,7@�t7��1�"��}Q�j��z����5�Qx��$��Tp�K^ań��J0��_�'ʑ~�A�j�8N�F�z�d��e�G�y�ȧ����HǌS*OZ�;�W\������"�vnTۥ�f1������=�� ܋��c�V��S�(-�2Y1�%a�/Mt���jl�JĘ?�|���J
S�e\3y�Q�,�TQ��K���@jq�=�����]��&v䒾����鞯�������8v}��P�[U�ߣ(�=">k��f�߂Ѫ2�͝����N������ݮrB`�/1Һϝ`��w���	�(K��5���h!����β�X�D�5φ#�푫�r�3Γ����>S��"
�P����`�n�[XJ�d�ݍ�Q�+�	>�8NF9�|��H�qMۅBX�:?�D����%U�V����V�Ǖ��T���Ow.��x�\�����-o"��ӎ��Np�"��h�/�mz�a�+��Ƙy�f9	��o0WR����c0�	BwV�$�]���V�*��m�=��~���|s�j�/aV���+�h�͂�R�w���w"���,�|�Z*�c������\K����Fy��yZ@1����]6GU)ڨ�!-�#�Մ/"��������?�����ZU�ܞk�P�?�hmח%�TN���7��1J��/,,��'⸾�KK{�!�/�vZb�����5s�@�W� �������C������g��w}�ϝ?O���IY��J�����/�,?wH�ym����{B��#�[δ�d��kM3�gΕ+W��xw}~��d�G())��\5��֋pL���p*;��9��Ɯ�,�7�Y���&C�lt��p���s]�X/��H�rS.�a����%���$	���@uD��T|5����gn��OC�׎U�jp�Oݭ�΂;D"����%zy��6���z}'���"l0�n�^���|L��	��o���R�܉΂�߱E�-�}�l��3G$�;�w{�݀��c[��K��b���ӥr���p��Oa%u����'{RRR�	�$��mwf�B��<�P���Ca�����au
���Ȑ�A�ڋ�i|f�P�ѵ�Ę����|����H��T@��E�{��jk;̽��E�D/R��H�b�xOk�w�|81ϋZD�Aj�� ѣ=7\_O�L�=�'�)l<?�wTC\N�:r�1��7�`{��ɓ'�[�����E���f��3�-[���bC�k�����	&�(�|ľ�3��O�$IzQZJ�@�-��Oii���!D$��W�G�����a��偺:RC����OpZ	 7�ؠ��H�Ș�؊O�=�~���	��(���"�j
�=m��|���+�
�϶�M"��	߁�d��$	)f��������S�q���i\�~��-�`�r��y��ڍ����].L���r�(k{{�&X;�#��`��-u�0r�X0(�N��������e�P�(����lœuTu��oAh�R�����f]z�L���$� ZG���U#�kݽ��=>=�l�5�L���f��/���D566�h��ބ�g"Q���=����ݣ��ޚ�����EN���jp�77���J���`�+a�@�m�3�������G���Eq���d5k��UH�<H��s�v6��|�S�-s�w�ퟥ:Gͮq�дLX+ru<^�#m|��s�	��75&*��;��[�=�o�kD�����ve�$�]ײ f���9�6)�U�^��e��U����Il�>������t$]ۣ3�bb%�Z"k&�?�2�����g��X*A7�	'D9��

bY_���)Y���%�� Yx_A|!��;�� !GwSJ����������D�Ae�e��@
�:9C?�)�ޖ��������.]�e�p�,,,h���َ�@��Q�h[*p>7����-�b{�g���Ucŉ�/kdtv��1���a(*��PfFZu�R}���A�d闓����U���!�=ؙ��E���v��3��a��q�0#�Y����?�$	v���g7h�ٓ�D�5|>_` ��d1&'��}m����H$R���Ç �|��
''';�-�7��F�^��K�Iutuu�2��L]`l�O����eH���G���ˋVy�zb����W���k
��O���Tuh�k��i����]y1r��g�s�E�JIH���)��?�jS5�Z%��M�g�52$��;�o�E*4�����Rw�rLLL� 4Wfz;::bhA�,�1Mob^��[����?�ژ�pSo	*zC(�Z�kq����@=Ka�ь4=�2�R�ޗۊ�o��	
rd��ױx
�z�9⼟*R+�Zx)q���o���}���I���PK   ��X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   ���X���5�  1�  /   images/a437e5bb-8d3f-4b3f-8093-72e2f97ca498.png��y<�}�>>*�,ݕl��d�=J�d	����-u�&�u�'{�ul�b,Y�!�1d��q?�������w����k��y�q�u]�����B���H���@�<�рW~;>��x=T�=��s����ϻ�zA _(?T��:�E���:n��~�6???!W'/+w!7O��9V�D��]���闉l��C㞲_��$⚟�	��eոI�OΆ{��w��y�V�Y��id&4K��ze�K�Ky�}�.ޣ�C k%��p7Y���:���x���T��"6��.��,��T^AXW��+���\��!y�Ϧ�U�
&S����6�h#}��c(����T�
Wsx��h6�c�B2W���k�w�Ht��_�Yx�Rǘ)��=������y�Y�	�!�k�\�?d��VS��(w���ؗ7g�usO��*��Y��Rc�О�\+�*Le����=>S�vײ����S!O9W1����@�k�EVS�J�Z���*��Ŗ�s�]��W ��ԻW�K�)�)�]�h��T=xϥu��}��j!�*'.�]�p�d���ic��:�k�|��E���c�#v�m��.����4g��~��t�I��D*��b�ѧ���kdU�"���M��6E:�ɰ��҃�s��k���PeQ\wH-{�Nv������+e �Z�ߕ����"���SfT[v�r�,_�I�޸�[L��_Xyz'�O��n}kgy��ɔ�r���.�]`0�*�f�xwV]uT1�t�"�pY0e�/ar�)��<����%�fy����[�s~��́e�D�q�fV@מּ/��&�'ېQ����i�\�	i/��x2.��O� 0���M.M̜�Y�̤]��G?9�B�ĭ)L��2~e�?�ƐA����ϸ̽{[�䶚(�RQƸ��^��^���&�@~�|"�>(Շ�tU��q��TIIK�uuu1
�ݚ?��Nn 9I�w��=��T�e��P�&ΆD��Y�j۾C�����M����GdN�d��<�I����~�!;�N)z��ͩ�8� |)�$;;� !��9_l?��F���2@��IĿ�W��*��-����2�pq3�7oor��Ͽ�w�b���	<�|Й��k+yo4~l�D N�+�����'s�������d��fy��72O(8z;�Y�e�c�S9jO�>~k-!�>x=�(��#��N}ROu����0�-��M�>�u<-R��`zn
�ɕ���"���ID(�0����v��伏���*r閦~�-���?ͭ�����ɺ�>��Kĸ�o@7�� �glC��u=	���/�����~�ڏeX�<ed�Ǟ�lwt��������g(��C)G�����ȦO���WφR����t�'�{��i�I1r���"�拽�5%F���?;�Z�[�;v?]�,�Ƶ
M2���擷{ڪJ���ɦ�GOKN�ev2��V[�,θ��[��`��%�,s��$�����m��e��KDX��9o��2[��
t��<�$cZ�j�#�����/���,�l���Z��4�(�
R(�/]V	8E`�dr�����:�N��Ν;����6e�'+����2,��ֹᎄ���F��E�\��{*�Pkfeî�'�ҍhc�Ё�K|������ʁ�ݫ��>)\�m����ӭ����rcj��N���/��9�98te�$z�j#r[.$W�X���O�&w�Z�A������Z՟�OѢ9	�ɑHEIۿ��"%,'�"˥��+�P����9�t����#|�w�JÉ��H���1˪bbbgn��.�SAŃ��\*ծr�,�I;�
���	4!s3)Ճ��������:B5!?4�Ɛ����e�z(���y)��k�ܸ�"��ar|w.����%�z_���j�#��pY���i�QC.,�;����{�&�k>�[⃈��
�e@ݫ�����Ζ͎Mb�2��e�����W+����~��z�m���/���5��1����_�s����㏚rw$��/�d ږN~z࢚�G�NOO;��Q&�����4��/g�����)�eC(Vg�PH���I�ӖN��,RI����ݎ�j��
b���/G�}+�[[۫���I*\�bb9EE���˹�*�x��� 5��>� ��*A��l�4dt����]��+rrrrdl�ΰ�2ݘΰN,a���̙b���ĹsS�r��~���G�鮩�`N |q	����]:'8\Fhu����/al؜�a-܌�� hשD<���X-�����GU����TRp�W��zL�������
�H�M��s⬣++�����Phih(UX����`��+/\.���Oϒ�?��`nE����k�ΜZ[[��W�mͼЧR�8R3�
�;�	��:k�E��6ԟT��@:�����	�[q?�����ev47W��ϑ nZ�0�1z!�at@>2��]��Ԍ���e���~�8��U�W5z.3�%/�&�F�/a5��FKڇ���e��}����ݕ�a��\�O�WF] �ڋ�l����D�M��6���"��~��V�v`�V*ɶ�@��?�P��V���\2�زL�nq7噣���~�� ֭�tnn�*g|MkT�J���+�Z�����q]�.kzvvv_��=���̡R��͞�"x����l`p��ቪ��5%̍��U����������5��g{7����4�8���E�_->tm"H��>WW���ˍ�Cw�GpE]���w��P�r�Ɵ��	V�F�y[m'����󎄽�G�SbYx!	�OB/�c�.�i�V���7����(�$������I5�� ��w�v��𳳫E�E�Ae�}����	x��Dt��\@���P=�A%��o����+�4�ɾp��t2G�
�I�rc?�鱨�����[���
�.���3��j�hv������/sj��������y�}��O5�9#�ݧ����>g��{��;J~�ִA~d��c%��hubw�l�(-�QXu6��=�0���R�8a.�)��Ш�>T�+����R3�;~4T�_扣�+�i�Ղ&�MI�R��E4M�E/z��͙�,xM_� �Z���B��}%O���j���Kr�sf�*)Sl1�z�JJJ2��U4$&�T[㄂F�~�� k�̛�b��ʄ��wc��No5|��i�M��2�x�'��?E�v�w��c�Hi������FC��_C��3�Ş$8�=؅N|��]P1]�n랏ۅ��)�+Q�>X�m�Ҙ�4������.sE��������>*"� ن�-SNmA���Ѐ��w��Aa<c6[�JI�?��U�DQDͯ��|��L�E{�F��#X�j����:^1L�h$�����N��\:��B�.+#�L~�M��쇹���G��B��!��[U#�Ug#@,��'������.J���k��F�Ƭ���ޣ[_ދ����PV�`��.�Hry�z =��+�ah��V(����4o2WWWqɻ|��:FnR�Kz��*2Y��V9�?k A#%��4_=49�0	�S� +����똮�7�퓃A;����C�I��ٯ]����m�6�2%�P�s\�#��S;Ԅ��o:݅ŧ�_k��:4%j�Tv�+9���7�^p[7R��m����{�d���%�ݓ��"��D�f���#OR�233#�@�)�x���ĺ����4�RϏ�����קꅭUR�h����E��]���)�����L��̛�o��x`��0��e���7}�[��� �C�lY�M)�����)�ؗ���Y����K���/�P��K������mԌah����S�^-(��1s�5��ԕS����]J$.N�uH~�n���T�z&�7L�^���2�Xݫe��kj�th�.ǡ�W�8ߛ�pqb���qÀP�m5:Ԏ׸P��F&�ի���`�o@������Tx�F���O���Q2����o�N衙�q�L)�����c淾o����E1
������!}���X{��m��� �K4����:��5e#��Å�.�V�0 �j�7�HƬL�K'�V�;�]*��#���m-Zaڒ�Zpu��CsQ] ��օ�cr���[m�s�u��A����56�u�<�!��cB���VO�u ��'жx�u["�Y6�o�L�o@�ͺﲒǸ^���D�ؙ�π�ey�[�!��*�;�8�W�l�}l}@a�����I&���O9.�Ҋ�:����O�"ꇻخ;�+rN����tF�׫M��Y�g��\�Oijy�q�G����`�5/����!�C�S'S!�3,��B������L��(-���w96��mP���m�-/��@��zy������<F{�0�!'�H�x鍥����5���w[�	�S-Az��6PJ�"Mqlt��&48�ܐ���F����L1�����6ވjK~o�hz�hXk�7���n�	�C1O@5�iH�fJW���;�~�Ϻ�W�Q�4��h�eKݡG��T��4i�B6�Ȩ� ���W�E��O���_�p�VUR���g(+nU�()^����ǩ=O���HJk�7<�2�7���/��@zր�2T��l���������*��4���lҨr�6M3ԛ���[x���ݣmw1#�5��;}�_�}���.��#��	�� ���:gCS���+�M���fd�<�U����9w�ˑ\W�;Ьjw�vX*��%��;��A�^�d��]�N��j�w؋��>�:?�~q�3�J@�g��bs��m�𶠲�|[>��gK�^tOtz=��nC�o��F��n�;����͂�

��6���ʧ6��3~Oo/tL��¿��?�}��ѳ{y'�#s����s��I���__�����mǧd��N�JN@�����kt�>�&QY�	�J���q83�Q��8$��l���q�,3-kp+n0Ű2��$�T��w6ss�/e`����"(�rL�ޞ��>��O��-%33x�'����u�'�ޯ�pmgq�cr�]�h!��I�w%��0�K�x��hp|Y�Q��b�VZ�~9�l�'H��,���+Ezvu���A@bs�LX6Xb��8��o����\�'�A�m�����9y�خ��o;��r�Nz�{w/�o��r���_�/�@
osn���o	l��m{��������.;�"c�: Q:;m���c^8�9EE}�ʪ;�{�Z����q-���ۭW/�=�|�s@b��N/�bo� ��_�\c@ �1~j�8�UG{�+�W�B���q/�2q�&!ッ�4�W�n��4)_�b[}K���
�!�|�qب]携�����I��dlkk+
���:� <������@��G�b�%��V�c9ʴ��Ou�C�=^�>�q�2-��!?@slq�^��0jay�]�M(B�&֪"$*t`�&�Ʀ���i»K(B�� ���R�́'�����=󯃯,�&��	��Y��X�=�������F?�u&�ʝ:]��Q�m�D
�����dee�V�) �W�6��\h��'׆*Φ�����=dw�s�knd��F[?���M����>>E��h	1����j��^ڈ�C.�.��ߡmo\������j�0�?�!�x�reV�`���Ͻ\Z�Iܵ�������W/��j�Ƞ&c�ߡċB&����@�4559qI�6��Y�#|(���C�Ҵ���H���I���jwCooo���M�w��S'#�?n=�LNN�u��\�E������sՈ��OLw��if�1I^�@i�L7�� ��^.g�ĩ,l~\���F���b��#��z%��,4s�b�8�Ք�(�c��ݬ�Z� ���C8�ם�1ʜ�\�CL�����4�7_�\&��LN�,GG'��A���m�J�\ �ـ����w�y��	�9u����?{:cVN:vqs;�R��^�l0��	�|!|������6k�}��b��\�yY[[�TZu��Zɩ4���骹a�ϭz�= ��vwNa�
,z�g�_`f����.�]��GB >]������I���ψy��Sa�i�Y��%����f��X˭��
ms�����Q`�� �Da�@/| ����Um��������c/�����ǯA "�7~9��m��$]<I�D?h�U <X�>)��>���Z�.z/sssR�J-NǛ��TX�u7�r9%g�H��^i����������Ҭ�)Ȭ4��c��(FY�r3Ӥ7�b��ڄ��^�3�`;�u����[Ho���(����ف�q��,+�aɨK�u�koW�F=��ӏ�������~�_����L=�˃���#".�O ������%j�s��ϩ�6,���xE��6u�U�@�ǧk�����L�O�S�EY��$,�I����8��S6���"���w.������'My�&��}���쭸�o^�!!%&��5���t�rf�7Zi?��~�̩e7\�4X��S�c�.��뵐I�{�L���@�u Q��`�O�r�VۂEM�����y%ۮXp�;#��	g��&��/Wy޴%��ɻ�,A�1RB����������<��X��R�?���/7�
@�/������s���ڠ=�7HHHH�����T8[�N�0�P�bqN7�(�MsmT�<������E�74�a�'+/_f/����,_!�,dDP'�L �\v3���݋�{��ak�_��]�KkRث��ɂ�u��I!�_�.�fی,�%n�W��f�t�������(}�Bi��^�
��z�ʕ���t	X���?(�L8t촆sx�6�[���p���gQ�������"�>>>��ɐW�����
$�������h[ڡ�0dDJf��<wf��+6��#o�������ʍw����ƨ��۸c!¥җ`t��9o���4eL�Zm�dQ
͐r�չ�/�?agg�(d|�1U�[i��8��0���VW�]k�HL�/X�<�031��O�"�4���Z�#LF�c-��Ɍ�g1A��p:W��E����}���
�k����Tq��<-_i26��&�%�?�:�U��#QL���7>p,C�֤Bv�=��!^�����H����#b�r�I �'��E��ښ�?��M�I�v�ڿM�@�N�)�����[�DB��YT��mLY�X}�R�zg����� xpp����wfo�=�K��ȫ��M�".��#`�^?��t�=��>7[���d>�Z�/����\�F��k��%�I�̜��T�����l�V�����CG�� �Z�-�V�����Vw�h-�z�BX��{�TG[[�A�=�WX���O���d$�����"3`�a��Tw�jx2D����A�er;1�B�W������j�j�����4i���h�H�`���ٔ�WG�-��~�e�)`���i������������6Ѝ��1;�CC��PK�p���稝~Y����H" }�A:;D�E���8Ĕ�`�n�we�r��*u[W%�e���6��χ�ɢ%��u���t15��Qfԭ10�k��c�򻩞��} �+� ɪ|�A�q�5A#�V��I�M�U,4 �hg�"�ѭ��{Y1���F`y��:&k.��so�N�&᳡g�����6K:`o}y] S�dJܶ-�)p{K�c������"����-c�@:��4�ukٷ�]_�3ݫ��� rr��B䡂W/P���1��7�fa����:��{��f����z OM�ю���Ke��O:��}�DY9X�#�8��5z�b�׹���F�@zlp-A�0�!�os��6��]�iFF���j���P	��ϵHڝ�w_�6��ƹ�A�%B@eZxznsr�����P�|�-��D��d���ә��)��p�����e��N�{�UL� =j�H�� ����I��Ƽ�����;�Y� WdSǞhR�J��ߕ����ЋC�� ������Z�:�5c>� �OUb7�6[XG�(6������n���$��6�����Q��9_�\�}ӯ��K��F�~O���l�[B�J�\VШF�Mʕ�:?�=�_<1�@��"g�rR!w�X�&A���!;��er���L��]}�'"-"��<,� ����S�h>,�R�TnBe�l�G���TCH�U\�O�!�m���ɔb34:�J4��zi�@:X�PgJ{_�f��Z��聼�d�7�Wm��.4���P}��u$mL/��� AP���g��,���)�A'{\���x�i\A�~����aVi�x�>���W��r����	��kȿ0��Ł�C���35��7��9���=
"�~M����[���b�O�qC�c Ĥɷ��џt.&#���=���[�!����!��6뉑?�w��:�b�4[�.G:'����OCo�*~{Ѳr�������&�q��e^���l���/�^��f��
.�{j�j�]���ͬ�s�w���7��sl��Lȅ-90�+�� :�ݳH,9�̠����̰Ok��J�g��-�	�ջ�Uj'��>�dCw��u�9���.��Ѿ�؍-f5\l-Lybf�HȐ����q-�N#ܙ'4�eת��=��Q���<����ʌ�%���3�&�p]�ר�t/��D`4 �EQl�:�+ah��T0,6�L�úuq���b
�7^�aֶM߻9k=:�G ��
����4�_�pqvg��Dn���n��� V�����w��zL. #q��n_�޴q�mQ������ n���_�&/��
�;�ZA�'���@�u�{�;1�~�փ��ա��͡<�c�l�S�M�����������D����l(�s����|���=u�~	�dh`�X�q`�}��r�������Oޙ ��jo�B�VỎ�&�/?��~�_��+�+��T8Z�4X?�*��oO��\�W�ڄb�yO�pɧ,˅0ˬé��rVєh�dI g1Q����E���Nw�ɴ��q�!�b���1�o({;=]�i�p/��@�����}5��K���)t�H�M���X�q�a=�W�k��*��R�c��&3�cRB�|���vz����� =�ȿù��(����'�I�sʅFp�J�"��;���n�?�Y&�2�4
F�:��@l;4��g����2����c1�������N�	:���~£�{��R~���"_ܸ$<�!���k*i#ccl̖�rQ�+R�<5?�j��S�J��Ɂ��nmlll���8W����b�3��̈�� ��$�����6���E׊�]�n�(��Z����*�u�VVV��9�<-�Xc�Q���hJ�^�9��P�MMuu��7��t,aã����zS�5\�S���
OI�`EiT�����8��n=����v˭��2-D�ȧ�-�lSm���;��Ƣ[�T�A���ձ��B)��K{��X���ho�x�U	�����1��T��L�"0�Ƥ���1�c��5���4�\����`YR��ꫲ�`�T���Lg��u{�ܾ}�Igg�|_|n�'���Mپjmwu�Xoh�I6x�+��l�q���'����~&�<���x������e�aU�Xଢ]�;)����t����={���°���[�T���*2���6��z�ӓ��Z�5���0��;�|�_��������ÃA~���F��)vs���P��û��E��@�s��Ff .�Yϥ�y�
|~�(ܰ�D␡r4���	'�+s��Z!!!�T�����Y�i&UV!�~/+w ���~M��X�?�VY�Ū���> p7Ӻ��g�h���^�*c�&�8�^�#�<�@(}���<�:8��qw���{����;����c���5Uk�zؕ�GK��h��q*�JJJ��b���Y�n�3��E���z��q>'���w/�8o�%�I��֔���c��؞������u���l�Ԗ�gq�"llY�L	�����8��ͤѻ[㯣����PE���,u�1�����
;�qײ��y�����k����k��Սmƛ�h�Y�V*ܭv���i�]�sق9�t�j�Տ�Ed=����ק����5kRL+(��c��#gf��`0\iG���̹)��}w''��Ѐ�;w��@��i�2�9k���� q�i�U�R���i��M�����z@��mw5`?wƹ���N�g�m1m9Ʃ�����#��=�L��3B�@ Z:����㯂ӓ,��I���ϝ��/Q3Q�P}�E�������3F4�)WR���)�b�T?h]�}'��,μ�|!�,��s�OZ0vr2*3$0pjoP����k���(�th�#�x��M]O�a���	Ĉv��@��U�E"�5�	�;�\��{��ϫ����*]�SX�� b	�7L]�}��|�옶6��ߊ��G&�nS��bBE۾��4�b`2��O�{�g�xRF��s��>d��/=\��Bt���������Kuyy�~�M#]���m�ֽ^��<�e�Z��G�k!z����X]�x����k�Z=���/o]:��;�����2�&,l�?���vX�[���$n����k ũ�ȣ�)�Ȯ�o���ozۍ?k���Mb+�z���~�ӧe7�ڠ�-����C��3�Anj����d�\�oۜ��������ex�J%�J��1Š�>-/b���P�BfWa�����k,��I_6�H�dm~���3��h:ؑ1����������]�o�l��Z���vL�ɌH�q���RI���jvt�Gb�UQ
:���r��j����@`��w����x������=�2������w0��ak�䯼H?��g:��1�.�ߏ ��H
��w��ι���q�Ʃ|�c��U_*���K��[�4&;q�q�Ht���8�E��e�~u�bޚR�tQ���,,!���(�T�����J��);��1uy��R�xw�tM���v��\.�	�۬1�2j1�9�!��uى��@�4
��|̴��c���m���"Ը.�ʺT4������5_׿N�=r* >�N�.Uo"�s���p�'�}Y$i�� �-P�z�Q�ɘw?��$��*p�:�=�V�X��˕�/�䂒v-���rF���E}�f��e=�.��2٬�5�۾�=i.�^����;�Y��*�ܝ�)�z+��N6�d*><���2/=��E��3��r��K�=���@C��sKEn�w<�@���|xv��B_wz�Аs)����~d+E��\c�NC$��Q�Ob9Fgg��}�5@���LQ.z-���=F���%�6@��.������' ���ħ���yղ림�]~TF|�uG��h�_���
�8fn�҈����<kϧI@�}���P��y]��G�<�Z7uo�U���ʩ5Q!��pj�s���;�]��]]���N�|nS�ͭ<P^Y��*0ЄG3sd�`|۱@:�<_��X,=ϑ�{Ӓڪj�|�z�����Qf�ｽ��.�/B�$!�໅������Ik#�Ad<LSA�o#]�`0ֶo�:�,P��7�'Tv)Q��9�x����^Ӳ�����,Pv�*Uݐ�LM�m=4v�6�_���z��Z��SV�N���K3��B �dB��zF.Μ!�rĦ�{�⟫܊c���m�(l��ˬ�R��y��_�U������1^x�`�3#ߞ
��K�Y��pg?�	��}��~�Q�1�8#BKyl�n�s�6�HͲ�̓�A���j�>Vb�����_�����mxD�p�ȿ�Lu�m�������Ͱ���e��}���a%]�Y����Y��ѧ����9��ˑO�vs�=Z7�btv÷c~˚�U����m�J'���=����?� �W�e�p����b�8s*t!Fj�G�G��&=b�&�S8z��t�Z\��@�ulku�N���^�K����:dܻ�;O�U�h��l��Vʀ��8�v��w��	��+.7�CCD��|yDj?�;��A�[�rx�<���	:�M�I�{��&����55_��$�,l{{���9D����a	cv�;)Qc���>��`���̳f���c�m�!}Z���r�����g���z^�tci�6m,��w�!��/|{�(��e��r`+ʴ.}��s[y#��|���\&=��{���a�1�j{���_h�74�^����mr�Kni�+h���J�X��'����>�ޥ0ĭy+�r=�4�i�{����E����T���?�6�'�3I�����.������=�Z���+����NE�s�Tt����Ѷ�W�k���#��t@�/K楣�TA��\�5�]��5'�T	_p�0������E��O_�-�2�{�O���xW������	�=r�Q��^�&��N��P�٨��`=�`����S
MGoձ�%�n1n�X�12��N_Ɏ�<�
r%My�~����r<�1M�X�Ǘ"�8p��1�__�ђ�����}vo ��^�q�LT����g��Mj�o��	��Hx|�/r���1�������Ze�:$RC�����`�|х�vnL�q&�I�\�w��,��=��~u]2����P��M��"�XV���@4)E#��uz�:v�
h�#�-����&�(�a��(i�1�3�t�hq��@YYbRy 7���np���1]�؇ǋ��|\]u �����	�,8Yi1��/���7����z"�Pc��j��X��.�~�8�!p���Mll�]���t)C�7����X��#���Zb�I�'kѢ�=�R3�Q�/���.]�����u�Gйq��bj@�c����o�xe�s��2D�Hӫ�P�f�%�d�����?���*K�����������yE���xdk��ƐC��(A�>�o!�(O3��"�X����s�ǌ��Q��X��ZF��9)靬u�����vk�ϟ	�Q����z���[�����,08Vj\:�k&?�r���a�Fò��o����y�i�k���h#��	~�222U�l�u��ճ�!��Kinw	8�8k�C�������~K���*�U��c�c�w��g�2��񭏟l�	rϟ
5���~beg{:�Q�V������aT(��t�^�[���	~� ���S~���]�9� �q�_@] �%i�*�O��]29-_��t�ׇ��]��x&�%Û>׆��dvY_�	�����Tt��+�U���v�e�]������&fR�Q������|q�iӶtt�>�C�Q��fi����!�����������:s|DrZ��0�YB�8a�$	u)��ֺ�����Z�X�3ۤ{ ��N�|�,iK�C�]��6�T���5�����D	��ѭ8ol������:~'�)����<ޔ�V���L~�]d�=�����X��	T���ݨ���v��a�'/��w79�m_K����17ooݜ�8��!nņ�9�铎�0ԅu�_״�*�N{�O+v`��@}�2�u�~�Lȿ��A��ԣrf:q�w[g ��̱i)�!A�
3[�O����w/fgy �BU�J��a�ࠟ4l�`j:$}���������G��ܧ��0m�������R��a�u�f .��n���mx>V�L3hM4��\F[�ӧO�6x-ۖڹ���=6�R�*�j�66����Ω�φ���jAS~?���Q.��Ւ��=������_�
�kE#X�l1�������T[�����ha��U!��;p�v+c3�N�e�N����}sl2h���g�����wz}��#'�Vt߭�=��.�̓X螁a�W��{��c�������=��d�tx6��� ��8TN�o4L-,�ZT�6-{�u.����u�ӱE	�.�H�����]/���<�x��͋�Jv�R�]�6���^O9�#�[���*��9Ga���ᕆ�{1�r��2��T5���B�^�������L���Ү9��vt쀻��`�CvK����#�:?\�?���x�N��{@��`�y@��f<�wTҝį�����w�Y.S�t��\�n�]�*I�!�!EDx�$��1�>�,fן{��`bT똔[�5�;"��،� t��.���HqyKj�L� �w���1X�:O��ƍ:����vY[?�!j�8��	/
�Z�wQ���h�߲����g�q����D��jLfg�_n��0[KO��-�82<�X�%V����8Tn��@Ny�5F�����O����|���x��"�0dmn�x�ʕ����"��p�A�Q����X>�#o}��
�k�hh7������75K�oP�X\�<K�拦ځw��f�����6
�'?Vm5X�,�g|��Ɔ06��.n*���Zf6��U)8�5F��E�,�9��l�EY��Pk�J\X m��������#�rӐ�x��z���'u�2���� �� �� �U����N���!��H^14S��:��3�}��'d2y�Z5�L�6����� ΃�����B�CP����c��𔑃��޶�; 3�Uҷw���k�C���rr&��W�
�r���d]Ȃ��vk��-�
6*oގ�🥚���ؠ��4555>�D��5��b�����!Y&`��a�{������ŷ ����B�ϲL͗t�I�(y�Mܱ�Y�{��﹠26O��5���Ay�!PN��Kxvlȟ�UaO��l��y��m;����M���e�װI��8���_p���5���?�TH���qCFk�"�ֵo4�b�H�j�����mo7Wn��z���2�}�}�F��:���r��c4k�*���h�����lׯ�d�f-����Nd8��%�A����Xu4����VUՏ���������r4`���M��1^0X�J����UaD�c��Ն]ݽs��]�f@��z���C�@e�zQo�p!�����
�y=���^���4��.���Ӝ*��t󎱻�# �:�2�Zw�H 3뀗���ZO���D������.�Υo2����^�yc��_Iy'S��{��j�9w���@)+j��D��M�Q�Ϲ���J#�S�^^�Ą�C�u(�]\��*��} ��pJ��������0��ժw�3��I+��ǳ��ë�6�/���bk2��(�w�Z�K�6�hjj;�y�.�}nʣw C� �Fk�~ʳ3���28@" ����2Y����Y��QyRڙ))�?���͠�;�� ޓo�ws8�>��˛?���-��Tm=;�����g�V�N� ��o��BT���UK�?P�v�0.	�z����7鉹��j�����P�J�=�=yC7˯��+���^ͷ�6�_R�����q�D�Ծ��JJCf�򏚿֦���]�8���u�GP�X0��+1������c�p��FF�ㅅ���$�7]� �6�r�c牧/2���Z��P��t?\6�띳�����ÿ)))M�8��~vEC�P�/���;�f�P������]�/;)N�W�E�Z�: ���oǮ�����y��:U�(�{�G#7�g9�w�o�)�v�m���c5}����b2ߜ8��{|��p�\����r����D��G���֯Ʃ|ۃ�|6\��a��UT��*\����_�m��i�R�^�M)Y�E�m?�r�h�}�=�@2�j~����Cݏ��KF�,x��"�0�jv�n��:�8vr�{�&�a�!�Q���筭�x��	P�qq������)q�~0$X�Т�����)�m���u��5.��O��zV�ֆ@��._ה�z����ӂ�1���ʇKGKˇbbb^-f����@[�m;��}y�r���5A�z�ŋt���%i7������!�RN�w(���悖 &�m�1��fì�HeZQ9^�i�zT�DN�J�:�gü �:�lȯ_6#���"r����������y�2��#�tNsu5�@@y6MGu�7z��3:����WR���>ܻ�Rg@��S�n����"�=�Ψ�6frrr���͚N��sc�4�'O(�G����ثb΀�°L��m�U��{�L���0�Jj^��6J9�}��Poz0.}���yP�צY�,�A{H%�\16���;��=�����t�X�L�u�BNmeO{��~�V�	z��}'���Ҳ��I*\ޫCy�w�M��.l�� ����>Ce暠���?�a-&��N��m�w� +�����8=,��t9�oЊ����<��b����[ILT��>T��-5��=�Zލyb�C��Yj��*g�9�w�����>�#/�L�ۣn�}�ǵ�鯿|�<��	:ժ�����N�a�����h렙\8!-���������޴L=�?��k{��՘`����*�\8E]��N�M��hI�I\Yp��S�U�7�1ŀ�^��z6<��
0���lL���09�\�`h?����ivy�t4�#��-}=��]����tF�dx��]d�`��S%�aJAF��~�o�+�S,���"�2��Z�/#.��i�b@a<>�n�*�pz � �*6YVF��2>|N�EE�������;h?�O5ܕD"ّ�22|��CҮ��NHH�Yqtw>�G�q �ذ�ϣ[�I���o�^�V+����ޛ��������υ��4@k�XZ�H�dF9�G_��L��fsk�M�x���Vͱ��AW�(K]>�m�<���u9JPP��A�E�S�MbD���L�|��͊uM�;�IG	����Q9��Ie��+�Ism��wWp�}%�2�x��7���A�ǀ��<Vq���;�6R���M�x�+W��W��X�n�7n��<�Z�_�`�� 	-�隨����/�&���V�?!<�{{k�Ʈ����$8,�3����[�З��U�R���M����A��9�<]��b�>3wy��|�G,x�UQ��Ҋ`2<C��ts�=�g�O��+&�k����My�t�ZS�c�Ԙ���H�,�֍��wu}\��
�<�9�c?8��x�N��Ud�W���^<����r�7�����XÀ�'�0�ص�0jW�y��9>���p(�d��>!������*���9 �����޶��L�-�����QH�����`�����>Xe����
�����	Q�RDI�P�%DZ��A�C�����n���!D�!%��;��}�7k�r-����}�~������n�ngf�SRRZ�avT�MG7�"�?�_���J!F�����~׫Q��֧³��e�Q&'���N!嚞N.d�l�m�Cy�[(���h��ִ�S����/�`
>tG�����S0'���v����;@kg���¡�W��%~9у������j����tu�菇Bӓᵒ���#+<�����g	ZVM�]�JDDD�� 7��^����<����+N���l����e���{��1]�#q�!�����g�"��6rBw�$ U��I���w~u����i���~����b�pgqͺ���9�BO�ָޘ
jS��Poџ�2�n3�ZE���Ɔ>�����g�}5*�2���]L\f�������#ex25^޹>H��C�>Qv��1#=]�t�<�~�5'��h~� �o��d�q��n�w:[�yoK�d�8+�9����e���a�;�۰����T��[Cf��/6��&�L9I��Ϣ����)�{�((A��B}q&���H>X�7�����nf}PO��W��m����^0,-ѯ`��X���ͧ�#��;�������󬓏���i��H�LήV46�>�t}�<�mk�ph[��[�Pi�{v�:�hk�v�h��D�G�g?G��;���s�riy�ՠ�ƽǻ4�o:��8��$�����wG�����d�h�+ZS����	fk��Wے�Z��&2�}� <<|o[���'nQT��ϳV��Px��r-2h�:�E�\�X��i/��ܗ�7�*��P�q�/,NKK+�9�3�n��O�q��2ŊD����gc�%6P���UWS�}_� �,�����6��g��`Jk��K��Ӏ���Y����:�3��<P�\Ec_Lk0^���֍�J'*)sU��+��uu�w%�VY�&(���Q�,�H�������FNx~����������G�Ĩj4KH���H𣐣���4���3��ZR��R�`��o��Gz�/gr�?w���(�}p��3N����V|�
dyHG\��S?	 bC�RKlA$����B���By
�읜�dV�[�7x�Z�'�ZSݾ���;n�	����rJ���l�܇\��ٖ�9��t��~��*�Ç��y�j�8�Y�L[(��Im�6tX����$a��ڒ'
�W�d����LM�׸�ţ����ty�.SS
�yS��)cri�=}����`�b�Qe�ܜ�NN7v<~�%f9�����RSS������.�i_M:"\�c�ż$��N�SE=yЯ�,hY_�����ayy�(z��d�.�YI�ޘKTW�`�R�5��Ċ�����Ф������ +kk��m��'w�
��?�?Ff�����dGs��p/;��f4��5T��-���g�/���dб�;j��̴K<�Χ��<�2�ž�:�Ӕ�!�U��!V$�tr7T7jPj������N�v�z5_m�{�ߝ���a0��~�g�fo����vT=�3}����p�Ս�G�gN����������S��&�����Ʊ���Rs����*�e��U�N���?�H���y���ǼӴ�"Q��<�y��@J�� ���kŪ��ď��+ͨ�ǉZZ��'wp�������K�W�-�,����&����Z_= ��=+��N�(�g�W�r��� S�]t�DHWh��p0�/�àq烙��<r��L�`.S��l�e�������~��X������+]���@J�S%�n��9��^���Te�d�Xuߧ%��<9D-C7�2V�|�R�	�7Չ����ƺ0��2qBm�K!ɚ���MƵt��T+�9X$�Z{.�2U9���b��6a�����w�:M{��g5q�h��Ɉ�kI?�ᐭ���J��y� ����xKK��6c��|v� �j�t�L��Ht�;V�}��=ٰ̼;`
�g����3��(bRRk�C]�l$�@�}��e�����5��߾ٜt����,'��89��K&��NFF6ʙ�m~EP�-�nR�Pcj]�����c���s��햖��G�^�����V��/Λ?I��Mbyo.��`ن&h�4ӝ̬oP����>�.��J_b���)��'���q����F�^+!q~�xD@�'}�N�{��q��q���Z �Ǵ�L�x��<���37�}���1�ʨ���R��Cx�� ���b�G�a��#ūR����127u��`y//Z�E@�������D=��R��dp����8��Y���bɵk�9�+>�t��B܀����]���=Ewxyߵ��$��~;�� �/�հ��k>�5<����=c[`����h�iB r��刣(M���l������4�u��[4c�\�����Sh�9�8��;cWg�r>�X@'!8/���z���08A>�}�'�Hqҁd���ۄݹ	��H�m^�����npn��G�����ߨk���ܼ�.�[��^�@T7�S�T�o�57/��9�h^�!�OtY��7��fη83]�R��YW�t���g��,;џ7�i�*'{3k�?�,��O�]��7vqF�C��K�k^�/�֪BA""~)A��hp�QH�3�!s�Ϲ�aU)α�W�ZZ�
I/{����ÒC������cz	����+.����?�'�ur���5��� ��*++)�0�ͱ�ٛ�:R�����(��_O3=ٟX�����
�PE��JA/u������Nm���{F�ӱNd�fzd��`������(|���`F�\ܗ�@o`A��"�Wc�����'0ҁ�d��bP�Y�d��&O�F.�t~(O�p^�IiJ��>�ce��RZKK�H���������ҁ�s|�]�Դz�����K�_�p��d����v���y4wZ4弛�a����u��H��DﴇE������B0���J-��i�Sm|E��E��EC�td�������.o�P��[����|�NBd	<>��Ť��_�����w�;(j�P��b�T���'�����K��r/�ή��Ti��`.G@��K�Pm4�7�����Yy��r��͎���-�; ��C�М���oHEOan�wt�]�n�������ޞ�(�T�+����j���j%(U�N�t�����|zEO�>�w�Ա*���@+N�k*Z�\�u-d}�M�O��Iȵ���cDk\�c�!!!�$-�QM���ͺ�fݲ@4|�VXh;vV���:�����h�r�A�_��>�c�/S������E<�����W*H$���ՕR��q�i�1��^�����>wq����2�6��Hi��� sA�-��o�i�|����x���X�ڵ��dWU�z�0���ӧ{�]~���� ��}HWe�-`�r�"h�I�m��E���@j��Lt��*���hC��3:B�gn�J���࿰���� as�qy��2���Ʀ�+K�$ڶ��y\�vk�h��LYx�?����L���e��VNlI*ϻT.�k�չ�X�~��)�~"��Q���!�����?t=��X�-�pV���U�2 ����tX�*��2��<�ֶlx���[q� �M{���{����	��٣?�����`5y�r�������;�j?��<�(,럙��>�k���������g+�F�@�s���@����i�5b/�Ve1WxTace�^���=��C�3mCS܏�$��hי-�D��;�vff���_9�9�I���LC�	Iע�N�2�!��S'����.��D�)E�pƹ�M�P	]0�?�TV4�i���Ⱦw�Eє?
��W���ev���L�);z�a������T��=�^���rmP��/b�d���X\UJ���Q��MP�^K�B���/�%���XMkU|�n9{!������)�W܃v$Y�~1��=C�8����]�o�����!���֔Nđx͡z�n|s��@e�����*��>Ӎ�o%3�N>�E���8J
k5�^��Xu���"m7F�ihp���;�V4����`��mv*o�����ʋ�4-�^��!P�C��=Y[���������g�}"D�Q7���9'�\Ӿϥabv����I킧_4Y�a�&�w��3�G�� v3�
��i]�/���O:yb�`�l߲�}�+N���TWW�PBI���<0��y|3;��B�V��9��[�1���t�_���RN	NO��<�2��1(u�l���܏��\Y��n�fƣ3�elb�H��>Hñ�Ib	�v�t�Gg~��$�Q��cccq�o%�)��$��%�]��Dc4�O]#xp%��7�fg�uj3��z����՘���-��	���d��ɚ�
E V@d����O�ӛ�6*2�Yn�)��ܿQn�Ay�0&Ӻ���x'�i�]q�w�(Xұ�(���$3��ޭ�ԁԺw�C�������F��QK�_��'�x���+]]2"�`�:e��g�ISVpx���G��t9ơ�I0��ǖ-̠�GJ(V��Y{��	�D�ǨJ�{���x̃7�Ē��{y�|D�x	�Xc�I(�`���Zce�ȵ� �/�NӅ4�+����Uȹ~w0
�3�tF|���s��~��������l֕X6�z������RG��JY�����O����������>~-7/oxv�c$Ϧ��9X��g��Rd�R�־�wV�YLz�-��ڈu��]�P��_��2M�{������l�5�M�c�Y�7��!@3OO��^Rj4�`O�1��v,X���������d�$���?nU�t�spX��a>�C�Wߢl���O��?�β��A�gw~��d�� ��9����uT��٨�2�ǩ��nX��F�*c��N���[�jg��_ڿ�;� ]6�?Hf�'ѣ�S�8-3�!t����j�ޮc����mL0db����iؒ?�tr��V{V&���-�9U��8�N�
�I�i�ɓv�k?ϴ� ��B�]�X�ۆEB���!��4��������W ��<өlsvB����x��'���I�՜�����cDC|�`���{��߂�Ju6�c徴/�^}2��յxѵ��otV�sh�TBz7},���i�%$�;����Kh��2�b�<���D�WUV�Y֢m�2`��gf<,?i�;4���E3 �֣�C4d��c�����"k)�=)�L���eR*F7ظT���p�Q��<�|��l�i� �?^��
.�κ��m��~f�w����c�":���E���{s�l9.]�;W��5'R��bv��{�CҨL%����2?��A�@�j@uۮ9��2�������h��57K<b`b9�Z}Uf�!D���KTzz�{���U��p��|�
�O j�>��`��`����f����-W�E�zq�S)�J�.�˩�ƶЏF�#�����or� R�c�]�)�t�\
�^��ǃ���O����~�-7����'wl
�p������v%�{Ic�W�	6+�z�%���,����˰ڵ�6V�?z��)Ò��M�m�7P2	�+����]JRR#FR��)�$7^��g�K'E�
��������#L��+�<>"��s������f\7�Z XB�p\��+��u�ӖC�}��qRL}�����*�y��aV�<��|cTc_1��3����1ȥ�OB~\����cU�ez���R1���Z͌�=�g:�^��=���F4I-+퐜��P�`|���M����T���k/�Gx����}X��0�͈�����6�|��Jo��U�y� >f�,�1cW�ݎ���j��E@��u{)���䢠{n�	:���۳5oqܕ����3:�F�w�8�S,ε�M�٪9�dr���
�|2ӹE�����/ȥ���`�������I�Kr�o�BYB�X�[��N�MnT1)5���^ �w6v��ˋ���	)AK�7�{���v�븧�k��'雺�hJ�d�d ����?�p0�;�-����8��[G�;�U�L�q�#�l|]f:!���͆����d3�{���*��E9$��{ׂAN��	��o�{j�X�]��b&o��s�@�	�x`���j-#�k�yy{�]�u<=|��j<%����茢ޙq�w#\�sb�}���z��� �1��͎��ؾ���丫�����ٗ��.��U=�ʚ݁� U٢hm�Gd�,8~ll
A%�����6��y,��hJ+ �n3��hX�ﴤ��I�D�s����t�G53<?��h�8����S����� 	W�a��Rj��������߷�QC�0J=Vu�E����řŧC}�2A��h���rQs0e�z�<q!�)�%�.�l��k۱1>��T�ےhΜ�fzA��M��9F옮 �LE�[p>���2�5�����D��D�;<��n@x%5]RO"&&v%�0����aٝ)�ҫ��@q�J�-y���y��;�f�J�ޑs�EE��N����q}����#��W���
$���g�j����Z(�!	�^@*F�[�!�Ǵ-����F���!ٔ$4�Ͻ������}�xY{��9}�����{GP�G;
م�:����-�,8�"D�ݭ��`f�Ieddc2ܻ��π� �~���}1��f��~���I:��S�)�&��z~��urH�7�WA^�������⻷}�~������"3���'XR�)�>Q�C*�SN����ԛ�]ZZ��vP۹��9��&�6P>N�#hJ-o�x���?����d��'�PKc��VNo���C�.�8����q�o��u���|��h{Z�\#O�U�'��{�G�y�p����[y�z�z�|�hG�]R6)�4_ͺ��,�4���u-�b�B�>��x�_�q�5:6Q��E[��p).��УEN���1M@�p���Zz�ٸED"�Y�+D�Ed���z�Y��D�3���L����p���'^���N]ߚ˯��9�+�4֣�}���S[.��h����p����z�G���B��--0||��1�����瞩�c:��t@����}}�(C#�E���3<�����.��Kc��8^�	��	f�dD$�5�M<��/�� �:Y� R#
��q�r���8�y�F���.8
5�-8uDP@;��G!!��ru*����4��z���b

X�HH����տӱlu�^�7�@����?��W�+hիq�^������"N�:+��}�=.��/Sj�/�æ�ҪoZ�R�~#��P�N����$F6L�,D#I�i��sݭ~U��j�<�|?���v�*��h���)x1X���%à�+я|���N��|�ĉC n��f�?���4E�q�>�W��7�P{WN��Hh��0z�7�
�)�噏��ke+m��c�_sa��C_�[M2n�ϳ]�qV���O)E`��d�}8[�"`߶ܟ�z-'���0���X ��|�F�����a���b	��AM�T44߫��6�L�v��K���O�o�� �]����;E���(-C_�����,�Ñ<�` �����V����P]��r���}�@��mc*��(,���971���}��Q-�hښլH 7���}h�]�^���(ٵ8�v"�m�vI8؈Ђ��;&M����P}-x��%5���q�e��3��5S�n>�R�_�d`��loI��O�$�Xz�Ϭ�P腍zL�̅�=�?�#�ek�fX|t_����tY|�?���;�n�𧗣�3�/���L����a3_�L8Vj��or{�Җ�m}B5V��~���;�~�i�E��J��/0��-��Ք�y7��i�����P�K�hu��
>�N�pM�����p\�	{v�ѥ]�1b!i�݁���l���ki>�m��oz�xUp����2���5v�$��<���/�ǊuCuj�olLc��#�b��0F^^w|}}{��F�u 0�P�.�K(���P>.�L�0�QA\=�H�yz��,Ab�c��Y>+z؎J�� ��z	22nG�l�M�8�xw�E$���u�(�>�?�5E0�u��!#K��h�Zws���Z�z�MQU��<�}�"�2l���,�r��:�ik"]�{;��(C����/�V ��hUV�PZբ��h�\�g^������v��g���Z^�RoQ�.�^�����{�
�a��&��OW�$v-��z� ��!
\L'{zP��'�{�v�kP����F�_�����Ѡ� b��5�p=:�+�{)s�˂5��;��,NZfP�6C��ݱL�{��q!�m����/44�nY�F��m�����pN�gW�ݼ5����Aj�(�D�F0�Th`Z��Q��Z#�p� �:��IaN��K��g�L�$�tw�C�f�]�-��{aKx�d���]�p���b��������iR=}O������qǝʔ㓯q��>�b�?�����n����>��˧����;B��o��{��8�j�4nu��>�����po�=�pq�c�1_oX�]�G�_yN����V�:��@���k��}1(�4{�B��޲��#�,F�M�N�w��<�^Ų7A���r��ݺ�>�˓��?NӅ�uwl�:I���
l/���WmC*[;�n1,e�O����I{0}3�����;�V��j�
�<I䈋~���y/����*��@�x\��2m��\�2m�C\&4��Bi��&e�8�I���=��Լ��Tc������1�9����� m�B�r;��:�3/�T$���!6_��o@j��Agޔ;�R
rr�lǊ�%���,�mj��قww�<����q�E`��)�pۓ���E�����x}#6���Z���2�Zi�\!�z�X��ߖe��p�;x���T�)OB������:�^΄�S�0$�IW����yt9�+ ����p���Tr?�,��m:Ӱ�]�����RR�c�Zmb��;Bv](^����y���5��7�*a�A����m	��I{���C@x-�ny�n��1.�ý��g�滙2���AvB
n1���KIZ�/b��-�̿���+�3�F��gUT��8Tg�������qF"u���˕jk�d����:��C���^s���p�M��5QV|���n\�4-�5�o�EXi��f"b����)�Į5>T2"�	[�f���%ᾩ��A>sM�E�R�KCCC�� �/]�51�,�互k�p��ǻR��;w�_���ar%XRG�_�����
���;X�oZ�8�������x㯅hjE�$��B�������-|q���"�Tk\�9G-.Dr��[�6Q�ٲ1�L�O� �1?�)-m<��Ѹ��[eeNPw$gUcN�ݿ'gC�PS��?����6�$��q� R����ԅ�tq]�3Ur������z���������!V�����+7K�}3���!���B��y*dv}x.���e)����ǀ]�l~�s�M{o�k.�\�W_�^74�q�}�2�{ute7-B&[&,��P��e� PZ���ճ'Jf|n�������������~DוD~S�:Ƴa��J9k��<'��x�K�U�q����iZU�p3�w�AP�� ��V����܅���~��1��qAR�`��ں�AEFp�E{�i��(�2�V�"�
�z��΁��X0`�V%A���֧>'�s�1%������>�j��_�Op���z�/C�y���� ?t��22��lv�;1k�=���5�"؆���sE�-l/��	J���B�Mm��B=h	_��-D]� �`��=y�����(^᪒�b�ڧr�=���"C!9圗u��f��SJNO�a�W��C"�c���	��u+��Y���GL�Q�.F�&9���F�;{�T�����+T��0�p����!K���H\�6�eu��?	톥�=�I�L{=��C�]>�FP��Z�^}���k��!�&%~�Z���'"���� �,�&��	a �u�����$�^�/ ���lek���F���&��[z�;(��Q��H��CǼ�d�h%C�u�]��F+�[@��R����6�f�:4�J�ZSgO�ҋ��>�"k�ػ�k�����L������|+���I�����666�[Ck�=�<h�������H��@H���}w�2�mq���\3�n�]k��	,��:��ZtB�Lv�V�	�}�u��v<h$��c�N������6�y"pH�� �{�ȡT��]x���I3�WW������i���[�Ϸ	��AMؖgwFGG��u�-����lDh*���)�B�7Z#����a��?]�Uz�J
�J,I�:L���3���	o��ܾ�2G���>�p������/?�>n �4댭�@-O\?�+<,�L��Tʅz��q%t�v��3�ϰD�sE�p=�._'���3�Nh9P�P��e��[���<<��w���v�7$'�oD L@ ~����9���>�w�r�4���h���,cL��HY �cWXiHڷ0��tv35d7o��=y"5:A����rv� ��WHU�d�E�
F���,g疢~�g�ڃ�^�>�>C>?:)�$)�,�����U��QɅ@���@����^������s�_��gk0�i@`���{�콃���Sw��`-ت0��Ď�|\��ϟm-�!ˬ��1��%�-�s'�4�?ӑ��l���
b��:3 �_Ϡ��~SK:����}\���ۥ�m�`e��A ��.nn��jir�ۿ?� �kYs˷����Pݎ���.�	���!$R-;�1��!�l����9��g=��RI#��'�ÖA���i :/�O>R�ż���4�]#g'� �4�g������=��U����Uڠy B�&���LCVW���������n��q^ĭ>����`�x^j�xVΞ]_O�jt�Ո~tx(�66P��
������1�`H��� ����Cr��*i4��5�!��i�ḃ�e���xucc0�+�؞�(���l*Zڴ�Y���5�6�~ۂ�H43U(������ �O�ٍG�a+����:])%��=�oUU-:�����߄��eZ=���5 ڌ'\��4��F&�k6�:<��L6a' �B4$!��7�^�O�J��ᆶ{GX$��T�Q5��AMRY2��p���+�z.�5^��[��^ؿ�����o���+�_��/إi�{e]����:�?��b����F�����#�wG��VLr��6�h�8�L�a�����	�l��� IuƟ_޴���ߍ��KE���4��s�˲c��}�Ĕ��H>E%��q�Bi���Y����g�o�_^�@w��4�:�Zk��KU��x�=���\�$ �zZ��m��"��+L��DĬt�j��{��e��.]����Ai�Z?�l��n��TG
�`/�&���N�z`���@sS�E�^6D��7%s*z��~�
��A�F����'w�?�g'�ryY�_��G�S��^co1�Mf�oE��� ����i�.oK��b���H�UB��m�J���`�]XX8/pi��w�>�ߨ�bƣ�8p�EZc�r+BQ��؈ܿ�"S��C�kvu������`ǁ�������H�Pi"���#|m@�S H<,��Q���"��0�^������ś�\���<���v����^��l��ɓ�6��QM��">"���/w�.3�og��xJI�I(�ё���iV_��L���T��(�u/�����m�5��X�S���v\��\�|�O4��#;~�S#s b ��/����������\ҪC ��~�8�w#�	��*_>�n/�Ʃ��ݪ��]�^}�+*j�b<�י��i}[I[|�n�uS�4��T�͋Z��w^��B�-������Oz�t���kk��M�����	IBq ���߿�@N���o*�f(>\��d"X��CCl�{�~�G9 �$5���������a-��h��y�`���0⺒�OOO/���nd���������`@'��&�`�(�*Z��߷���<;�{�+�s�l�tЖ�e-�բ"���*nA%Pbj�υ�אH$T�h�]z��� ��(Dc^I{�z��gf�[za��Z��:W�:|�����s��s΅(�ٖ�����'�d�Q(�1�պ��aU9��z��|��!V������ة�DHh�0���f�owH�{��ctl*l���^EF�27"��f�15��,j�T�����FC�ҷi�������Qr	��^�z�B�R�Q�
6M�b��\��M��H��V3}��F�Ȉ��ܞ�=��{�r�A�ny��;��Z��þ�u��slŃXf�ފ�{L�K@ ���)ZT#����U|~ݬ���|��̤�P�w4L&�p��?E`���oE)��WQ�:��l�7iln��B�I�/Vx������u��DUIt|B����KN'޼��4g��Q�!GMZ	�Sj��������/f�K���mx���@K�)�L���Ka�������~��Wc�h�'<�xK�g�ְ=�Y(��0�bY'��$ �5
5�:uoJ���W��f'��ґ�t����aw���o���ob��6'M��,{���nkS�/�&/�٩r�h9c��ԛ�4}i����/+�	��g9�
ǖ�o�sY���������C���^���� @w�q��풏c���r�E�ħ���F�[�б#�ylT�� TJX����}�m��=�� �Ӄa�}�ωKe������APA%��*���r;��dg�}�A�IG�Zx<w��j��wq2���|�n�#�C ��@�v��	3�������}NT[J�(ƅa�hIr�x,�iG<I���&	�g	�1�����5h�9�ڠx�#����/�����{6A��I62R���%�rÙ5�r�+>���i���a>�v�b|��s<٨�[ы�0�����v˃`v���#N=���F����waL 8	M�m��@ �>�����箸�X߾}3+.D�d3�qPn�,F�$=db��<��T��W�O�6�b��cN�+�:��%{\29�u�?��m�|)�C�e3[��C�P�}�]���9�{/3cfb}rd���4lҒ�|�3O�Q����O?� 1�8i��#\�HƄ�n�?�z
�y@��6�Q�p(TW'�,\�������s�����,�gįp��'췞sRSS����A?�ᱜd	�����A�wI%+�`N΀�Ls��Y�Jc/C��u�j���g��g�{|�.�-�Ywf��?�&�H]�c��dP��2�y+���+�|�	2�U����T���-s?�4M��s�F��V��
���W[B{w���zR
Jf���TOG���e����#�v�7΃b���%�(������?�@c�l]�o���UÆ=����V�^�9����J R�t@�e��yEYtDm킞M�D��:W����#�L@�mo�H2���yZ��l��v�	��&JwO�}��> W��aqS�'�c����&��3�3���{	��q󒀚é�b$g�>��=d�*�I����3g��lj�,�8��k}gy0#�n�6�+-�t:S��۱���,���v�F[[]���g��#�~+�ƁA�v��p'�����~�?���|\��vz��D�  ��z[/^!3'o�g�4((��h)qxj*�c fJAj6� U��<.�5?�[;h(���n�q�z�R�qď<1��`v�ubf8��i�+}@�u�G��r����[�<@V{�	�`��#�+�|�����`l�)Zi^��ϛ=�(>ȣ�8Iz�$%���O陮�n�)���#rgE������3Q����� �޶/4x�`}..&�#I�%�>�����6����t1��'u���VR?���l
��Z쟤��ڟXG���׿�f�������ZVv6ε[�-��ė����@q�.gq�.��e�,�:��>P�.�7��sj��QG�8�Z�4 ��S�$ OR���] [�s@�N�!Wp�s�#���O�s�D����X�8���rd���N��Edj5^��ht��[ *F�d8�# �C�sm���;�����{o�!U��!�03�eNK=.��s�׭���#Q��\gKN�[ކ@�����w6�myϝ��M�<�q���g�v�}��<t�G�t��X�L�/��r��`ޫ�=��Ts��C��Y^�9�(L��� b߀�b�7�HP���!�U4Q!G�ä��l�C����wC������K-�X�ed��K��1�+6��X,�6�����{���X�\�24��3:;��ؾ�O@�-$v����KM/��/r�W%ظ��ST�V@��e��1`��"�O8�,�4�� �Cc��ٲ��y_
nm����1G��"��2_��w�s���)[�0��� *a
�`����C�����#=��ծ�:6$�n��%���O�K�%������C�Vh}�׎�]�n+��pn#��%�� �U(����&�95d˜@^��̊
^x�늑�s?����s�'��%�OW$�[�֬�^���3��������V����Ff�����U�v3I}����u��;�9�@�g�Jf� ���Ҽ�X��~Z *u�a�[�S_�6�ޠa-��\f:@L��R��	Yȿ~3(pUh�Pr�+ �HxR�zD��u?UE~3�I�F��"� ,����q��쩨�v�����vo����l�[��0�c��9��쪧c��/���$�*ٓM ����� �{�+,�Ǌt>�������}OYC}���N4��� �]  ����;�����m+@[0�kyev�<Яt��c3��@����s1���"��	��N'D[E/�ˑ��Y��e�}Q{D3i,�&��}�61*"I$��6�OA��Rw�[je�	�(	*"|�ϫ�<K�,��3a���C4��*�~w�|̜l-+EM"���ȏ����:W6���ν0W /)@�@�(����\m��AO`z�{��I1�� b��5Ӆ����Nj�FDD��������rj5�!�d�}c*��Ӿ��T�c�����dWp���� ���MKNƆA��� 6�J'	��%�AS���eGL�=�2{�d��	1�ܼ<���� 젿�EU_�ˌ�(&�}p�+>�K���:��M��u�<�MM��A&�?����ݨ��������,�yK�>�,�b�*�����b�"'��5�ɣ�͡�ݠ�*������Lw��9���"h��;u,%F�e�Gd�C]	M�'�.<t�-]��ί<L?z��鹓Y�vږSis��^-V�TQ�Ũzzxv��+�'��1Ӝ�Z�޶Ɖۻ'��7�_~�f���ꎺ}�t>�`��E��y9Cù7���G�.k��؜?��QKX����E �g�����1������$y����z擩�bg���������#�m�F�g�������O���	�ic�iT�R��Y/����E�E[Ó;�4�إ㑛��Y'Ц���ם�k0��;?{I�����p��]\���|F*�ֈ+��D������6!J��>�V�����OZ�7N\��|n:���>��*�y����d�^�bߤ2� �n�	� C͕�w����������wX�ej��	I�x��m�[���
�`�˩B����AB;�T����.��]SB~�_�&:n���@c놛)0Ԯ�<:u�������9�=�~�	4՝;P9$�n����+�[��_�� �%Hh��I(ğ�����R��X������x�����/Ǽ?��!X�� ��̼'�=�����jK�����y~- �y��N��f�v,�$�l��@���G �c���K�I1xVg��&RkǼ{w7I�LL��uC������j��$�`�����JZ�Pn���ӝ�j��h��qc++f1Ó�l�X��!J�����Z�G��,��rs�J
�2|���uh�KH��e�ǎ	�o���rI<�Ӗ\|4=�</�7����zUq$�&��d�����I�i�/�,�QM�T���4�h������V*�+��^^^�9�­"�5���Z@P�+}j���u",ŀ%��^!g�Q�g�RP�B�8ZZW7ő����Ǉ�� 3`��1X-n@Rs��qVGi�����9h�7
�C �''u����z����(Ҙ��`���X&P"�Nr涺v� J!Űӌ���q�-��sj0T������Ek�D� i_s���2�ŧtj:*d�G�6T~b��Q���?gՒI��V#.�������L��8�*M�e���~�B9�2m��W ajYKɭCm�E=��!�\|}��8
%V���(%9Y����X\����)��V��7�HȦ]��ff��x���eC���;P@��|\\���#� ���$>�[�/~���=}g�P��h�}P�t�˱T���Gۂ:�
ia1�S�0�(	��g��1f�P޳`$�+��U�Ҥ	`Q�B��V�@Cb
���ݍ�����eE}|3���a �NN7�=�$�>��	G�ړ��|�2�+P��6��җK��2��C[�?^�)$I���p��X�,�q��E�J��`�"lC�#��K�Q�����s��r�B9�[�<}Q��cr)��[���L(�^X���e���������`�x�98`�~�F���&9j��������+�U8M�Jk���M�O�k������K\q	��"RN�7�q����ry��>�(g�1�<l,EE���@ .�X3�'r�.˳$O
h��m�I����z�8HBq8�e�yqv�J�̓��8��y���F3��x���'f�誐�l������M¶���E���.���깜$���ԘH�?X�w+�x8K�\)\�5�f��R��º�z�e�`$�J���`]	T��UH~�����mh�Y�C�"8vK�͛7/����{��Z��Ƒ(5馔�3h_)~�AJ�Ԟ��W6�o\5=_���<'���z�_e�
�>
 ш�v���e ]�%I=�J�ԙ*�� ��QK��`���L�)c��}���#0�gϞ���}hw��E��e�z4�>lVPT�T����<���d��}���5j��'u���
Hx���B !fJm��=���/YQ�Rm�%�6 t:&&�58�apԏ��:,T�U3��r�1}���>G�w��,��m&Ů�ӒQX���뿱Ġ`w���N�����F.�9��jD�� u�3�;�&Q#!@��T���tM)�$7��Tz�zTh9݉�(���>�J��ț���IA����:���P��n�>#X;��Ȉ�_��;�i�i^n��cCA�u��"�1��~�����xM%3<:������C%�c4o���9�K!�,g��+�`���&�:[P�^���||��$4B8$P�:��c!8bξx�}���y�H��<�� +D�yx(d�@�٫Zda4���P�$�r'J�_���.�qT��'���/�	�KN����$�٫r���V��)�Z������ؤH��,Z$$#r���n�%���rw�V��DZ����D�Ĵ�l�L��bB����g����|��s>���<������w��s��~��v)UA���X�#���fQ_E��C��n &��m窘'����g�yJu
�:2��sT��8���9έ2Lb;����̝�~�>�gTK����XB(^��N��WC������I��y�7��������w�^hXx}P��O��O�J�R�Tfn����/.�9r�MR<��q����ۜ*��8������:�x9���!
⍿�_'vumhA�N�������:?�~|_C�!�pg��j)5uL\X�I���\X��U4��b�cc�-�� ��9�R���FR����?���O�L�� ����M����ӻ��,{=8�2�L�AJC7wE�B:rhY;�Z�~Ȅ�*��m؎��t ��-��DW���R��C�Σ�?�>����'Ƞ��h�{���F@Bݗ�2a�����6'~�ę@81::
>������C� �`X1n�����f1Ƹк����t�]�kH��{����U�[�������{Q�4q��4�
��`�Ğ�08#j$'|A%+	������<o���/�� |��� 4�����^Q��p�Dۛ���D��'{5��۳Q4g�6}Лm�}�S����/=�#��։��,*����?�8�*pFH|]j����/�1�A�{�2�0�$�-B��r�L�#�+N<x����t�%��|���N���tJ�Jc�n�ɚ}��f�NDg�,�R_���A싿`�_a}Y^�r��S�F^bwb����/�C}��%�{!?{z�= #	u��Ŭ�䏻N�ћ�8���ȗ�y��sו�{I�VBv/�.˘U������_?�h�}!�����?u��Ԗ(/m!�}��ұ��N�o�NO�^����؍�Y-�YK킓n���DE����t�����?W�X����Oߘ=z��m�I�p��I@�N����m���b��0N�ݔ�R����Қ�eͰ�i�C\n��Gs��L����ٱ��)�����N�����?��@���p�� ��t2�v�9;δ�|M�YOIh�,�e�S���vDV�_}M���1V��|�Bu���;�q��kS��ZsZv�'x�ui� ��T��m��� �U�������M���`��'o�s�Բ�Z�c~
�qw7-C�1p��;ځU��wʁ�am�{,�Za>�wxm�}�S�T�ۭK�y���Z�%��5gv=,��11ۼ��cEi�3-&Bы���6�¶paa�,����Ͻ���,N����&���@���$GK�єX^Ĕ0PvL�e_�k��<��C�x �^�J�<&��I��ݗ�x�g���0��i�=u�W?z��G/G�t��:Ůd/BW�v<�g�f_�5 ��:�(wʗVO1��M��-��[���q*Ԛ�(J��H�0oE2�k9��hn�DW�.�g��u���Q���6��2ls�]`X�[׀t8}Oؤ�z�Ʀ|n�`G�Lwp#V�N��E��Ս-=>)��W� �d�0�.X� �a� �v�Ttk8jI�&)�a��WH��ݰ�n)����Vm1�����g��{ya�sn�@N⩧�����K�- ����͍��?"���y_Z�@O�NM%>y;�zVP�;�[��l�A�V*�u@K�]�\��<�̞�P#� 侪���2
�V��勪�ϕ��P��Q�����'~l-5���o��!��5$+ ����y��V�5])�a�3$8���^�/���P>�#B��w����h��ZW�LI=\#�nO�㈛ۚӓ�d��ٛd��7/7��oQ*1�{ -������\���ȩ��?���_��K���cuC��Vr��^�D�Bcu;�qq�)��G���� ����Er;����� z9�R����J���WՒB;+".~[S�|Iuss��:��b�C��S�F*��N	��5����ֱ��؛xf��c�`!,uu������A�EQ�	�<
e�i�L�jCtce$ѭXe>�-- R�������-�N �2l{U�Hy9N[\\,!��'��Ù��`0�����W��gX�Y�S�1A�usí�A�m��p(L����?��gef֟���V+v����j}t �.D�ܜo�8���e�Q�r%�~C/;.�JZ��9�>�nU��1�cQ�1���F:��A���J�UŐ��������9eG�v�Q�� ���2��g����v�j�--�7�q�JpI�
���
׭���)�i~����6����$���p��Ļq�0%V���%�g�����#�P8Yfܱ�@d��cͤ������355��~̖�J�<�H�5���7C����G��WX6xvWUta)D�����wH&UBo��m
��\0h��]x@D�F�_��5@�"#-s=���yDN�at8�뷔��!8 �cqa(�EF]�5Pj�3���(JMb�k���3��[�P�KSqP��/�J�쵥�|*�ߤm���1�%����::��}�e�	�!���ȯ1��m���T�Ǥ�\o�b��"l�<<??_1����PC�a^D����Ӫ�+�rz�������ZW����(#kE��ܯ�g���,m�(�=���������%z$R��E�͌,�/���/PK   ��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ��X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   ��X+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK   ��X����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK   ��{Xw�'<�  �  /   images/bef45656-42b5-4670-a699-453aaa19c38e.png�YeTг�%�nda	�E��kI��^b%��K�������.i�F:������9g�3�a��7w��U��qipQPP�d4�I�?����w�U��8.
n((H��0�o��?%5\V��l��p�F����9ٻYY�Xs9��f�Ҡ��~T�����:21�B����l�1*�(WH���bZQ#�,Q�Q���C��T��DA������I��׃q�t�}��1X���PRj$�km@���1qd�j9r��YG��]�~�Y���WX�z=[��5ҵ�� �G�2Ǧ&��PI�c ��p2���*t���7F���3�7!���X �R�Q�n���aI�2v�̩���A����99��}�w�ܦ;9�l>`�E��8�������Yz��a��O��W�q��O����:3(a�{4
�u��Wᵋ&̪���F<{�j��kr���[���mUY��KR�x�P?�%�^T�H�m�^����?�`�D���Fm��H�w�⡂s��&L��B;�Ґ��oԒc�MR\���������![����Mb�'�o^u��O0��'� LP7���9X{^�=��c��m�(SL�clv=���п�-o�I���QRּXI�)��A2�v�����?�jj��G"�Z�\.gۻ�)F}{��J��� RΥ��b�zL(�;1.��>	���Y����^��cD>�A"��f����Sz]w�m��a����8cAeE�ʽ��8�+0��Q�
A��*2�<Q�b0Rz8�$5�9ˣ�U����t��/a���F�$���>��ăU��VD��aa�}>	v��
E��幫������m%���iW�:��	o=�{m��ڜ��X�z��T(�^�xPG1�36WA�h^����aqly���RY�?�����Q�1�LFv/(]��|=��jg��X��\V#s1π��ļ�*�D�]v�o:��K�<h�^�Ә��nO�[��
�X���Ɏ4pc�8K�S�p�[���*�>�;$	j#C�0�'�,I��3gIi��F�U�E�k]wS/c]p�ܜn�:P��8�cn�0�_�ު�T�1�Sa���)ۻG8�,:�e�PQ�ƛ�Pd�:q����B����U{`u�g�`�Oq>29�h�6����%��9�4HO���7�(�_%)#U'b�GY�O�:�9�W�ܥ�7��,�]	��S
�2l��|��z���]���^��^��Xß3����f>�(M�r�|�5�K�&`�|�v���Vz�Ԫ�^m�y^�
��U;�&�����&�U�S�'jϧd��=�ڔřQEh�%�Zfp*q�TTg�`͂��K.]��ǭQ����1���䦭|��&�Y�o�HĈ2�$�ѽ�嘅*�<MJI89���9�ֿˏ�X��͗5�������Q���Pl����}Fn����Y�w����雅&�|*�V��ee\������#`K�7���di�/@�H�ᶗc����� �2f�qp vug��>�V��u$�*H����Қɕ�����n]��5��*�Lb@*~�Q�Ah� V��9`�j{��
��@N<4���p��*0�r�y�J۰�1� �Ef�pZ�4d�f�5�L��F/�V�@�z�.�SLeC1a�H�ڍ�B�������~���ݠ|A�� L�Tx'l*��GG�]�!�3}��+Ղ�[����<�s�<w��4�-F���"w�J�\\�!����Js��x�;�t��e����O^�皈����w�f�d��/8β	{ύ�IXh<Aͧ]�"��[՘��Y��n�?�c��ގ'�����$Q���k�u��J'z�5����'\�/��}M��[!����@��my�w�v,�d8��t���zrH!J��/�8�9ɯ�smdN��<وD�a+E��x�0���8f�����c_����n:c}��4�``b�z�
���b�D�P���L���@j�R��k��q-�O[:?�)��+�MD)����tG�X㾕�D�]��2ڟ�*)�Z�dxy۾���(v4==�,���o[�T���QbE`TfD1�Lfm�p��8��/{;��Ze�u�s4~���ī�������uO��cno��o�OX˙,p"�m~��496lNRU-��go�`�[�G�j��3�az�|1��6 1����t��M�+���s���Sh��5�?O�~'�v!L�n�p|�c���@��ޠԟ�g��P��7�aY��]��"�P���[f_���7H�\'�2�y������pM��d�v��NKѾ���<��$��6E��#�|o�t�7������v�?�N�򕋑)������(��̑�{�K��V������1bM~$�ل�*A+6=�͑u���6@gN�ԑ!��g�"����Nh��b�4��r�5#P�>���g�4�ӛ�q�ַ/B�z�a`o�6<J��*�mt��"6����N���ö_��|q��/g�1��M��l���5f�n�Vs14X�,,�l��F·����S��})�v������Ppy�X�:�N�E����%��&/�i�l�����؝>�~��{�=W]㉞a;2S�1x�G�y�M��|���U6�-�H���]��ơ4<+v4�ae�1e'Z8�Ύ����~ȿ�3M6&��t���$k��
K{tg�X�l��o�!Fd��Ż$	6丌iho��7�����cO�P����J %炏�{ 6��Z����dSk�W�qO|�:U�̇�	�߹N:g<�JO�g�e߁�{��Jݦ��UBD�'������T�������䆘,aI*է���^��Cn�<� Oj��;Қ���bU���/����WE�t�M[aam�����޴QY�v�ɧ��8|~�L��6kI�&�|��݄��ز
�[����4�l�۸��9/o���Q&�ox,bOK!:�ՔzX<c��IB`	����Ѧk�q�����N�|�Ƕ�]|����4�����jx�=���G�݇��_ϐHU'���j|��Sdot>n��Zg7Wl�룳@��n��`.wR�vA�gwRs�m���
�E���~��2UDMjH�2:x�Cӵ����*�9���E����dɐC�S�K,66d�!�1���Xp�qS�#��8����1!^�,�̞�)��+�0GX�`Do��[�w�k���*�Ŀ�v�����o��*��7�R�-���v��gj��e��#Q!~��?yxW����}�����&��֪����CA�U�%O��F���-�E��a���K��Ծi�q�uS�f���G�h>�*�1i���
C��L��&����zz��O�+�/�]}p��m<<�XfRX��'j)QL�3��	������:^tű�q�*�PQ�I�0^B��l"pp@P���,��-Y�죷$�7+���Î���a��SЉ�vb\7���a�#f�.N���e�G��L]��$7��Z�m���2���Y����Xf��^��2�hT���(��O�)�%ԊL��W>,
��&��dm�{�ew�>��� ��e������ǅ�m�qF����{f:���l2�$�vf"kb�C�`&;`%�����"��:��c
by��C��g�����´<�]��~2�o{ ]�/�(u��<*��~ �e5��D��6�ng��}�~�p�D� ��+Z��N�f�>b�F(qGg*շ���s�$n��5/�������Z� ����҉�ٜ¥2���1�E�����pW��,��ߠ���n���[�p�Mx>��f���xd���$P�a�q��Y��{�#���M����oi@LnU�U�b)��՘��_lm��q00tX�z��JU�6��[c8��\r�U}{�y6�awp�P�Q9���eCe�F
xD K&Q�'}!TϦg�����2��o������ٚT�u�G��ő��/"�2�5�F�e2�,Ww4b��e��k-K��7,�BM-s5�/�&d�Kͧ7�\��c���ù��v
�޺�iI�.��Z3��E-'���_����'ٔU���*�� 3�{��!�
��w�L��X��
Ņ�!8xO>]�ԛ@��_o�=<0���%������P�ph�H[��]k�9�:'X��r��l(N�J�l���AQ�Jd�qjQ���YT	�M>��>V'Ts?ܫ�\T�s�H�Ǻ��"vʛ) ibF,�1}�NR ��c�}I�L�C�Z�P��P�MR-?=�qP ʕM��*P�����}5��TG'�9�J��ᐒ��ˢq}V��6܇蓜�C�aT&5��2��Ut���-�#�8�m�؛�)
�|zMP^ݤ�;�+���ZI}�������)�u�,�3{��{uE���6^���p����d'�	n�X�e�~Y�GT�b4y���y��4�@D�e�6b��%����r[hH��7�����4J�67�D� �;���� 
�G�xBm��z�o����8�vp�s^���U�"���!}�%KL��c)d��YЄ�����6�.?G9|��0� ���f���ޜ���u)��ڤ��G,U�:n�T��@4Ck�.��b��#��D
��EA�s�s%(��B6G�s��o�x$�!�!�*eO)Y��N�٧`⛉(>��W�F ��A����M��G�f�+�J��ƥl)~~�g��J2C	vh�n�?0���Y�Z�㢾r��?�5]Ei)�0`1{����u3��O�xF;|xE3��a�w�t�7)!"�R��`x[P�^�]������"2�v��Vd�"���=����i���'<��MQ�Lh�11��Hb8fc�3D�j�,UM��1$�f #�t��1��>��P��|�oZp�����|����Z��@&����\^����j����F��a�+N��aq��%jm�Pt���p,��@���)�)�ʳ��戟6���I�s[s"�E�t=쁮7�{��X_����1������O��I#���k�W!�^���
#�j�c&�Qq�I�ʳP}��C3e~�dZ��E���}LH��	�΃��O`�j��*�MA�߿��"�r�I�CzS�~Y6M�
�7�J����n�*�Y""�3�L��K;�V�(����M{+����)Z�%�Jy�ȣ����T�M��{�ai3�Ǵ"今K�^@����V��(�����/�-@�5���5�a���CD&#�'Zkn��Ԓ�jf�z(�E���o�wH��=�RJ^��������V�9�h�7^Znt7�"/����F�6�o)WlH�*���Vx�3���%>l�W_�@Y��$8N���e�Sw21E52��g]/v�	hy����c$�9{�r-4�7���[zw��:7��7/�c��,e=9L���Eyx���{��ũY�H|h/�
��0]f�(��|�PX;�����zU���w�%�}<IZ��d��0�;�me�z� ��/��̈�2,�n�3����ǟ�ا��:}�E��a��1��*���������,*���cĦ�ȋ�ʩ3������S�T_�l�p=*�UjY�J<SI���p��yZ�5�����W{|�\	✡�o��i����>6�����a�W{��UB�H�C�i�� 0�Eg҆�rԼtf�h�V3	���P ��?����0�D�#V%��0����~@���R���ՠ��b�v����w-|���Y�l�D�@i;� �C�;W�T��c-��H�&Aެ���6[�f*��}�Tj�7/K�S��~������yI@�<�^*�y3���8ա�^�r�\s�w�z�I���&��T2�ۓ����7�����2��`�=^�X�&a'�^��𼓻S�p��/�n��v���ˠT��H�qi��#�l�ŝ��ܰ8��X.gr]i\����E�~��z|���	����l}
N�	����Ki����V���u�hV���^�wv�	����~sCM���
cb.�����"���(����n�ޢ2Ck��l0��5��Bt*n-I��CFR��9�i`���C���,f@��'�C�̲= ��į1�$���Aπ�(�y`��OJdD�q���zO�b�Ot���,��=�-��EO�޹1��qa)�򞑧�)w���ٍI1O�d�##����rcǑy�u$�6����)퍭:F�5��и�|�=��8�դ�^�~�К�!%�IZ�$ �ز�W���52��sm��fx�#.MKw<�ǓwT66����0E\�k2w�r�$%{�p�B|������b�>9��i�nI��j]�K�}0ߍU���[�yTήzM=�y='�� `�ӕI	u`�r*�[�R�I����ߟ|)@Eirx��4 �я39¡ۻ6�.((2�;Ȣ�3kO_~��i�:��e��u<��u��b1���+��V�$�hUh�gB%�B��ߙ��ǧ�6�}4$Y�9j{1*��m��c�@���&��,��u˱K(tqbV(�6��������Υ|���]r��[Wtaq��Z�d��ی� ��9�U��N��,����uy��-���ȸ�����E@5_?b��A��'��eun����}��;� M%�9��k���z�:�h+�̟�w+�-��t]vh��UN}�X�f��P����Xn��UZ�M/�F��fn���9G8Y��PЋK�]�G�oւ~�8;e,�=�>�Y-����3�l�/Q��Y��I0K�mL8�ķ��W�{��^��L�A��&���u��k�:V�k�@	s��2�-�hm�rO�Zܺ�q1�=��`�HkL������=�D￫�#nk��f�7?�ͤ�|���/��6Z ��g�y�1
�ތ���J�_����u���Υe�T�Q|x~�ՙvm���})����H������qڑ,(r��Y�Q�R�>�lrϋ`Sg�}��Z���+���o���ׯ9B��V��2;|=�|���m����0��7��V��d~��]�)��V�˥�0��/4�e�BF�� 3o���C�~��'&�����������=Oѹ�_���<�h�xh9w���A/ٿ�ޚȟ��7�)���ş��G}P(qt-���uB9#�-3i"V_c�"�S�V��%�C�)�����J�V쀵Þ�Є2�If��Qt��]Hn|0��e��r�c��#���5I�L�����Tn�)[�o��]Ჲ��f�X��)b�3q��T�#~��[�*T~�1���=n)7R������ë->�R3>5��(�*S%m�?PK   ���X��g)�
  �
  /   images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.png�
!��PNG

   IHDR   d   B   �s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  
kIDATx��\�k���߻��d�dK�jA4F�H\BK��N?p[���/�C�P(n�R�?Ч�ҧ��o�@����UR�QS0�cl�.�lY�W���jwgz~�=������������;s�~��9�s�LBD�O�<�D�B�0#�R)�L&E�\��j�*����$bϞ=b�޽?��o�YLNNv���#dvvV,..�l6{ƶ���,�;*��!L
�{t|�ɓ'o���v���#d߾}��ݻ �;��n��������W�92H��I�z��h7"G�Ç�����HR^V�h���e?Iȫt~���Gt�#�l� �aQ�>�����C��m6�����F?�jK�Eİ�~�O�^����/؏���m��\.W&���������!���bbb�P>�o�V�#D���������
gΜ333�T*}�:��'��h�u��3���=I���b��	D��X,b���v!�o�p��
>pR���={&8Б�G�8u����ܿ��D��d)�N���3�������;�������"GM[1�] ��1��$ #.;�|�����z����N�:ձ�G��+W�xvg�1�T�P�����uk꣏���?�޸q�#m�!Q�sB��	�2D�uP�7a����;�B���MY��۷E�!�<��!��aw^y�uw��!��:>�!�t���'�����ѥ�·��"�Dx��dv����y�cc��4.=�����vD�t(��[YY���L:$ ����d��w���&����(��P[4g~��='d���.ҹW��&�v >YU�&�رc"N����0��r�:�P��ᡡ��r�cI"J�&vtx=ச���?9��[u��r�DMOOSL� cy �H�S͝0
�F����ˁ�V'����>H�#�0Hm�I$(��. �	��ras j��J�!���_��x0�u%5�OJ�*"0!���h���������d�C'.-/c��*O�m�ȧN�C$�.��:�UҖlo���˷b��ϋ�J�a�	�H�(��!��m^�0����͂���P�\I��!0!��8#T��`��ُ�2�F@����יt��,����BH�������>̕4��k�@�jnb����ٞ�(��5���`�7
�)!L4�
��2�'�G���SL 0!<;	�Ӹ�L�I���	�t�2Sf�~eɝ�a��`uez󃖄@l��4��4! :�7��,��U�&�B����4��.B�d�I�m����u����*�ج�;o��@�����J��.�v@�=��>h��@+�v�����κ�iG�:.!~e��< ��?M�t��ۅB[��݃��&o��|>��:jbB]uBM����9��J��!rX�"š��;�{����G��6U144$����V1�׮]���T�g	Q��TWu���ctl__�$!��q�������c/^������!6�����t��9}	�"��t��gGVΓ�;$%����~R}������{cjjꗃ��� �7M�����oY��3�.�:nCԭ��N�w��Mˉ������$=��e�))�f�I��`��X�G��g"�W�.]�300�aGgY~����_Y��� ǹ��s���]�X^��xNrT�K��xK�V�U���1~�lB�y~�h��Ż���;`�k\7�Ћ�Pw���z;�M���8-T�JKH3R��dB�`9-Bt��mZiK�XH���u��#=he����K~�/�-�D�W./���4�W$;>�m�����x�r@R5�|n���!����!��U����9�V�??�mC�H��u��W��Z�F˄�$��i���v��V;�����*�<���cx��6&��sq���"F�P��':�`?��OB�#BxB 8��<[Ӳ!��� OL�#�-�	���dI�+�I��ȟ��6ꬲ�V+��2	Yu�/Gk���5�!�kE�C�:�WiYe�yΕ6��D6��m�0G����=�>��C(���5ǳ�Q	Q��F]U���!->Hû�ePG㍫?Y��5;��S	e��T櫵r��)�#B��$�S�����E+���)���-is��CTP�Z��~�����6|ޟI�*"	��B_��7)��ׯN�<�/����9�8j�!�mB�0��Fj�-L�Q��8z�lI!vw�w�f`qH����fg��ŭr�r�5 �~��Y1���������+u \k����u�a2!��N�:�\�{�m�N)�D<�X®�˗/�x���m%>�QZ*�ga"{�&�JHPpI

+�Lf�}�K����و ]!!rX�$���Q3ݽ���9����SHR�I��%�7Kk��d�jB�3!�&��u��&�p�~�\i��E;�ʌL��l�I������#5C��l�oT
��m\;�]�����׌j1M��BB,� �
��8n��{���!�n&��Hㄔ�ٯݲ7^v�Tn�qJJf��,�?	��{6M�]��u3NȾ�����<!j5���%���p�-�M��m�	+�z�R�,��	I���<dD ĉ���P�\+���:�nW���t	1�.�T�R9�n�B}	q���|������۵bص*�
���7K�X=v}��P	�?l��v�l��k0xO�n�����Wㆰ�v    IEND�B`�PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ���XXs�銙 � /   images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngl�T�m�6<Cw�t�Hݠ�(�(�H�H�HK�tww*#Hw)=4���>�s�k��Z,��c�s���M���2>5  �WUQ� З  �\,�'�~��oh.r�����/�E8�gl' �������.�C*WE}W]GKW����l]>�;}�u�l��� �
��=3�=<���1���/�U�Qq��hZ���DĊ2d��s>�u>EYẼ�SP����L�H:���pt� ;�y�o���P(C ���ȁ��e�$���)Й%vݚ �������f< �٭�=���:*�������0J��	���� Ԙ *@F��u��}$�)IzFf�Y�	��$��;��8d�+9������%F��-լ�u���{إk�o]s���W[�Zx��d�Y�9��$����ʹ��R����a�%燷[�2S������x�9�w;2z6,���2���� H���m�z�#�2"(���	�X�w� �/�q�լi<hk��.��\�X��$O�߉��s�g(�4'eh�j�w����Pښ�ᣔ��'�K�sI�NY7?ι�X^��2����D����/�<2��|�|���F��i�ŅƮ����5�H�Y+u�7	з\��NC�/�����dJ���:�^� z71���'"��gl�n$�n;{��h�t����u��va�"��bEie*�S�c�#m�t${F�滬�k�уQ�9��v��@�MW&~�[��l��Kl7��v�^ݧC�>-x5����n���,��XQ,�����Od:/z�γ��Z���Ol[��k�c�,.&�� �U��"���mކW�L�x0
�����w���MZ��P�0��-R) U2o�Ng�����dt40�R�r<�:��qݦ��L�,%]�+�ä��SvxA�mc��}��O�C�Φ�U�$�b>3�\t4 (gn���'`{�'7|�K��h
`h�F��[Q$*��4����@����d���55�y���=��$��n��NmgD�85f����!oc���_ز� 9L��)�)��1��G������ڈ�x�N��m�0e��/�-Ħ��T1ɝ˟p^"���� ²hHF.>M�<�n��C�#�d��YT������sۅSV�Zx�������fwD�ԼX�n������4z9���|�����e�2�hC�~L��c��Z�¢}�Ο�7o%�ð绡�p��}�v�=3�M���� v3o@�R��:�i�'^"������e)��u�����_�J2��R�d8��'�s:*�U[kj���_h>��gr����͛<K�>sN1	H�=0Y�r���{����$�^e`�E��"d4,�S	?��� x>{�_;�˚ě��������X�J��T2A�@�'�K�P$��Y���e�R�l�MR�$R�㺪B= ���o��EZ��8K��`�$�40���Cˊ@1\�Y�ӿ���'��-��e�Y{����Cv�:�m�V��o����mj��Ԑh>qz�'!j(�KO����gn4��JyC3�M��?��"��`��M}\����{�\{t\S.j�3Sst�߫��/�8T���3G����6�gj6����O�0�=�EЏP�A�v�#I�����>�����e�|��}�N	��¿���#��+ ��RY������/��W���K��\,����u�>�u�mUx�N��&�n���K�*ޙ{�L�e]]�˹���M���Jюt�+��^<y_e�<�[2{�8����@��AbZ�k٠<�:��V\����A������/�5EGg1c}	��=���%��~�ߍR��p�f/i~"�T�>�O��:�� tw��f�A/9�۽�d3K�X����mh
���_aߒ���;��^��˻1$~ZJ���}�rz�=p�e��w��/q��)�G��ބ��[�u��](�l��g��w^�8���tA��I
je���R,.t#�o�b+��ڔ�7����u��H<�I'�g�����(��Z~Nv�5��h]�1F�R�Ç�pw�$sC�6$K��q������t�ܭ��:Uq�-�AQ����?Ni5E��|�o�ڭ�5 �Ǩɿ睳���3ﵠ��� �ݓ��Aj�s�>��t�v;��\�����;�d��J֮�����P�8�-�{���Yz�OMGi��Z�������O�'�{�Ute�P@b��fO�C̷y�8c@���:�������M�G�X���6dտk\E�j����l�dʛʴ�/e@��0����o��8N��
���]x�)���5���!p~�i����-3���Р/8�r����>}m�#�4�1��A܍	;�0�-�M��a���%�� G�<����6��`ȏ5مt��u�WtF��{vhb�Ѝ10�h��	��A0� F,����4r�@;�Z��"ŎI�]�[e6�ޟ.�.�v�v����x}R<�_�)2���Ǒ~���ms!"�(>p��:g;������(��E�n*�����c�ͽ�k�mD���3Z��&��s^���p�e��d^�36,�sl[��S�8��U�+��_����EC������?r�٫�3�Lf��,m41��[��@��a��偳�/T�N���H0�F��v�6��8_�)"c�J+H�ǋ�;�u��@XƣF���������������i��$�ͧ.�<E��FbH��Y�t#�I��C����XJ�Ya�a60��p�:��޾�B���Ft�G�\��~_q��4�~�_Y�rt�/�D�8$��Y&d(�e��)z�po�sqA���/w"���/,�ܝrWC[X|8�����9p�LT�������O��7_�8��vd7�����~zN��+���E!�V�F��_���r��m�m{_&�z����˄�F�7;��+t��i��K��
�>`Xei^K������'N�Yh�W�D�&"��ٌ��yQ4%� �G$�K�?�yw}G9h	d1e�����-�<�:n0�x�;?���@������\ڶ�~B���l7���[A��ޫ'��g��љU~�B��㭊Ac~x����z���,ɼ	D�%m��廓��j"�x;X��|��4������]q�{fY'��;�,h��fe{�[��(!����L�b�=EϬ��δȏ��۫G@�Ԙ4�KJ=�9n<ߵ���hu\��uG;�d�/]�-�)W��NqB�E����d�]Ha#�?J��c�F��zZ ?�]���c,���VL"zlO�1*�&~mMݫK9Qw����S�K뎿�_I~r�g�c���m��)z��D�6֝������M�b�0���.�q�5�ܑ_��O5�>𩫅�'o"kE�]�q|�u׾����s��"3Wz���Dv�#N��G&qz/څ�U���P -+�k#���7=���Omݚ���%X�m̭��`�f[��̋�X�#|�!�������j�H:�j� ���$��9���2����l�8�#{VQ���$����I�Id:ȊI�.��)�����?����d30Naպ� �C�
���;:p,��׫�$`�13������SL��׈�j��[�Ƶ���wz���y/~X,�2v%Ae�[s�=�Bs�ܦQ�7�f�v�w�
���p=ח�N$b��+`ǹ��B2�;�،�ƛᲱ2S⋢����S�[�%���T�d����0�װo����>��}�b�w�t���4��F��kw��@�Ad�}�<��cmΖ�seʈ��O�w�\ľn����%eR��KLli� �5�C0	k5L�����I� �����A��i,茽YS|<�,L����e�hX��Tx�.�Rqd:��ғ��t��4�E����K
���ʀ���
b����AF.v��FV� ��Ewz}j�i��T�sz2Q��,c�QEY�e������lG�E}%���Oz� ��!���$_C���Q���ǃ�O��r?����1��6��W����u؇��L�����;u��zco69\h=���1)��}}�!�\׺m�28s�fVes����RNb+��>R����U�ǉ��'�4~ :*	*ޚ�+gϥ���S~v�$��-�Z?��O^�{�,��B]��@JC�����(�:�ެ�/V4-~�`I��9��c��
���ײ����X�k@� �m��q{&]�
�����Lp��_�KJ8�9�)tc�Ke�ےϔkl� �w&���d�UZ��I|��)H0Q��A��Zry>���ˊ˽�y1H���|�T�g�<����[�Xe�>mC���~�~ؕ��sz�������E+56Џ#\���L�X�>��d���o���/����E@Q��Wid�-� qt�n�y��+����X.mԚ��yҲ�d��l��B���]S"�&? }�䑑�M�޵�^��ؖwU�e,���h>b�?\�!���Ҍ��e���N1mqz^b�J��.��+D'j��(����n�(�O�[��;W�}����r��А�+����U��xI����������Q��9��[_�[�x����RUi���./��^��N��1=��~��;(݅Y�:Etl���(���� �̠1 �|$<80$K]j�ݰ6|`��x��L�)	o�td�<��P�{5OA�g��ݜ��72�,>�H�2Gz�x��k�2C+�/7�`��|�^p�fvڕ�l�3bVr���<]m�ø�W� ~GNV��z�#���"��LΜZ����1&gI��O���L~�j[��c.�e?�
��kMS��G�)�<e6နO�V�W���C�D��qL��E���ic��䯗����{�n>������˕H?�
��	�/�	�̽���3�i���:8{<��B[m9���=&YI�,�B��iz��<�=	���X�l����� �	�f8��1Dߔ�zޥ8M��T͔��tߤ������Kk�o��i��䳸���r���l?`� �5|��G�y#���*�i>ɒ�?}�'�N���2���֙���I����γ�兛dmB���ӟ�c��f-�<����'�[d�fzX��|B�����ϙw5�@v�c�~u�z�c��L�F�~�rd2\���d}��"�����9:}�I/w���)���L� �0@5c���z�.yϟ�c3od�N嫮��u�d=d6�囗��a�v����!�w�ܞ�)1s�u1�2�Ѥ��@�id�T�6�%i�Ef���ﴞ�U_d�k.��>Q$rz���gؽ��S�SQ���u��>��.6��1WvsKnsK9!��dZ�_��/e��$�wC�|��
�(��y�f�e9ܲ.:��l[�V��~�㸄V�IH�vvn��[~�/S���jyСl �jf��y�2>(�=�����&H\��%���{��t��	=�8��G֝�WP0?����/ ���o����d����ߋ9��\:��7�c�H^6x@�!;[?���v|�RC��1��R�& k�S�ud/�'3m����($U�L�'�Yh�����lCx�xƛ�֐���Q&\��U��TG�!-�5i���X��O��o<�B�u-�%�O:�C(�S��v�"{���͗���B݃W��W�)��?{���!��u5���>��7��dG]�r)b!+�AQ��>3q��VO����2!cPϕFv2�즪Ө(p���ӂ;v��/���S+�����J��?�0�Qj�u��xF�Q�R�c����HA:|�u�J�u����'Qe��7Ue�;"D�nL�f~4�M�5�1��l���2CX0��ݰb����E_�l��9��L��A˰��k�� �Ar����uzG�ӳ5��aQ 2��/t�j��5p�LF�i��YD�;�N
 �5chŏ�x>G'�hQ�9�L��uK�u���&���Y�t��[�f,J�M|�X��S�)9�;߄ĦD���C�Ԡ����a��y[�%��v���*�p)W�D�f�Q���a.XM4ף���{D�O@"V���Q;���������}��^��ɪO��hf)�gG��_��Nۋ�%��+��Tq�;?�c��'.��т~-��W��T�05)OpYփt�
L^��\�\mw�@���'k�Y���8�߄�Ғpy��A�R��*G�|M�h`�,�l5<����	�	h��/�Kr��"��A'�W������x���$N^,��0���؝�i����Xr�w=���*���Or[s��{�>;tI���E0��?�7��9j�R�p�)O=�f�U^�B&,��D°]w���O�tz�/�AoE�=<��d�%������+�Zд4����~�Q;I��
"�DM,�����أf������p�U�+�/\�L�^q���eGY���N��/qh�cKHwmC2%']�L�:0�Fe��f9��	 �&t���0o	�����)tZ�4�K�]�<���K�t���	c���߬�3F��K�(�<��%�bՖ�#J�齷%�@*���>�� ��#$�􆼝��&%���1���)&i��Z��`+w5��:ݍ���*f��ѿ�d�|?3,Ji�b���<^T����p�ņk��0�|����ۡ��܋S�W�>}>�y��+���v�#Ba�h�0��,�0�q��)�[�l���Dis$�)$>��7|�o*�X���?|9Gf?W]�ovmmJ��'ZW�HJ�bC�xٶ��\ \cNU<t�L���Z:ª���+��6k���v	�j�[����� K*5�`���	h�U7��S��]���1�o /���6kf��U9�J�;��Ӣ� o��`�>���4Ma�hd�`�_���2���\�Z�����ϸ���*^�]?lӎ��$�-�h��R�u�H�r����� ������bv�?�WU-�nV���d���w�T5�\JH���]XL徂����('��5ֈ�z���jjK�Y����Cr�����V1�rE����|)mR��4�m!	W����j{Z Bui(5w��lg���5뺂V~����8���k����#�ꜻUGe�U ��=}���+�U��q�`l��)��k���r�g4�ŕ��M��N�����5�E�1-�	%H0���'��Ƴ�A�{�9�C�����nf�,���cm2U��yI���c
.�T������7��F��R��3�u˪�d�h��ڋ�υ%Ju��}$S���D�	�&���,286X�5#G�q�>4)?{Q��.�ۋЎ8
�	>����:�] �̬�q�owZ�:�u��-�m݈8��� ������D�ñ��Ñz]i��l�"�[��?������k$��S׾���:�k"�
��w����& 	"T��
��۔�$T�h4/15�Z�Q���Fl�K��!An��ݷP~6���TPp�E9�W[ـVT�F��'|(��n��3ռL�e��}��짢�Ds��SK&��m��(�	t�j:ۦ"��.�m��aU�x�d�\��^.�����_�w�ӓ�dS�g/Cj`���_LB�:�m�F3�pd�M�C�����i��o>�Db��J��d�+B4N
��]&�;�ߠ�1C������z��.���l*3\���'8h�Ǒ)A���l)T��E0mT�᳑���;e���5:����N껫Wo�Yr}�����s9\6�>dj�T�xfd��^�=9��;��[��x��ONQ���E�3i�k�x�9�l���[e��O�4hl�e�_�QST�҄�����+�"�2n�j�F᎑�$��T��j���e�Q�"�H��wl����~so ���+����4׏�:���ʦ+�缬2k� d�M Bm�,�ΦMq��a��W��}B���BkM�;����;x��B_�㻢�>u��D�7�������ז�`Rk�H-)R��y�#N��	;sUFt�ө�6�$��Ƙ(X�葚�@����[����Y$m��Z�oK9?^�lgdOk� ǂ�
7?2StF4�[���n�pv����Ҷa�с�y�q#R+�)6�t+k>x�ѧ��ϰ�zQ���h8�55�sf1Qvk�v8�K�D�%�%!�.�G���|�HO,'����o��k�1��Ntdj�c�2@QY��S���^d��5�AH���a)W:/3�������P����=D����PK�G��CF��J�yk.��f��a�N�>�<H��(�z��8�!��M��vD���4Ř�Q6��Ӹ�	 (ԏ�Ea���������s	��"Ζ����!9N�q���)@���T����l]��i�;����u׹�K����ƺ]�>��7���e��^6�,ҷm]{
w��(�[���J2`���A>,����-%Rd}��.�G����QSP�R\�Ʀ}��E���y�)��)�ζ����֩����D~vO�[G�m7���<���a���H1���������q��������佌0�rdP�`m����c�e�O-����b��:�x�o]��C��ĻDs�$\Z+T��ij��;J=#F(����+%�(Mtej����o�U���e���"�%6q�C�F��q�L�__ѳ�y,[�o C~b�O��b��q��5̤��B���1:ZU�����|Ij�1&��xlj樝f��y\k��Ñ$�ʄ$��XQA}���گh��3��_����D��!h{h�zYO��l_����9P��m\�R0�F�y@�.!_.�k=]j��>8%�%�,]Ğ� ���+/Σ���̜�5����r��uL��r ��7Sc��:��0~T�p,L4�r�еSW�b�S�=#���Mô-��D�}�eؽy{@in����F������|��W��@TG�j�ͭ�9}܉���q�<�8����`�?X~-�q��U����%�D�39+�x��Rb��-^�:>�������;
"PყK!˻ER�5M)�r���l<�YD��w����p݁OZ).��A���S��s�D�Ɋ��ЁK!�␍*O-���s�{Ƚ����w�s0�s�kB�!&pfh����I'A%�1Z2�Or�\�]��j4�j�������-y%�%�o�K�b�H�}7\,��7����̡�M*F8������>�fM	y3]��'�zry9ǎ��sP���ђ�#�<��A���J�N��'Th����Wna������s���jѽ������9�))����l6�/!�m2D�mM��f�%F�d�#�O��ZoE�WQ;q\BP���u�t���)����l�z�7�ެ�)/-�s� �^�hH �����6�h�W�\Tյ~HS6��Y�ktl)��1l�z�������I�E�h~�5���殜;�;����i�衴3;�r�`υa�1 ��R���$A�[�%e}�fMQ)՝���hǉ۽��t��B���[�t�x/��
�����u�y��d� XU�n���H��S_,>jۥ|�?>@/������խg`�F�8�dy�2���_�bd��Q*2�xn:ۢ�d:���|�ޥ��L|��R1C9���9���;B}�l-.0�y������q�/d#�ц���4��o0���Tr��'B�����~2Nt�=1�[�a�Ù�bCx�[,>�M�lٱA67���,���oxĞ/����Db}��}�;����,}=u�_Q<`��|h���?����^r�3'���'����W��d#��o��
�}�`�,5D#��`�u����2�)9��SͧW��*���sJ�!�0sɈ���#Պ�1<6�]�
�I�p��0-EJ>kF=�f�;}��EaZK�����׀f�ʞ�8�_���'�hY��c.Ð��8�w���6~XUg��}(�I��#����r����c�fvM�Ͱi,�S��l�PH��������ټ�,�X�3|��D$��8��7��T�-��yBb�/"C�?�W�+f��T	�����T�0˻�^�1]S����`�Uf���l��a�w��+M�>!�g�e_nG���B*��H�G���d�>��/muZ�/�K��/
�̒�b O�y�[��,W�rkX��uT�B���S�.t�ĭ�3^5ݟB��@��J� S ���UM��7W������6�;aT?~@l8U�odK|�����! M/]�����^��u�~V��M�Gp%���}�����|�(�GTsJ��٩-�nV#����Ա����	�*�E�]Fng��"Œ�p�⮌Z0�C�V�qAj�Z|8d��viRSf�+;�r�������a�8i%��i)�qf&��H t�P����TL�$j��m�ޜ��w��Hf|Q46�V�f!5(뼕��c'nl�V���$^�`�^'�]���ۖ�X?'�W�E���q�[���-EtV�q	����J�H��/b�,v�p����3��=�!����hi�VU�4Ŵ��A��۹\��ɲ�F�E �+��06�C��#�H�1���up��p��L��|FaM�}�+�S�����,5Z�������="��ň�"��~K1[��9j�c䠥���i�Q�a��<_�7ft�8,�|�5~��њ���g�h�F>YvI���ѡ�왅�&����#�	�1j����J�xn��������-�=��J����=A�P�;�p�u)e�5Z�[�`���@�Ծ?��H��/��Fg�}��.�MM����{��?d����&�D;AF���o���^j_���e�$��Bs�띩
SA* /�e9b�J�P�����ԚY��iT�]n����|ᥦ$�d���?.�4\��M�PsE�
��E�(Q6���aE,�������u����`yd�
���e��7
�c�`��>a@x9$*L��_��w"��i�sؓ�஫�@�]��+�p�|A��'���Ռ�8aHfX`���|�H�W��/��n.{&cX��]�X�`�N\k��vB(K�D��I�ģ�n�"�zeͭ�A͖E�k9�We��d\���7�%uh`�dp`�}����k���Ԅ�X��/�U��~0�m�z�E���'��Lϛi.�O��S��t�w��J[=;ks#pSi1�����Q[�^! $8��������+�/*��ʼ�Vu��H��U�F�gK��軠5���5,]����}T:���+��%_���;��-�n~_���WO����^���j�1&R�G��#�.W	 W�YdQ��)�[�c��&��B��|M��*RO ���1��#��y��l�j�e;Y����%v�@������w��!�	�hc���d9�+m�-�TW�x�zkR���E΢j�5(U�5�|i�DOy³q��6�QID�v�6꒿�h��!�M�T�,���l����*��sd��_��X�bJ�ٝ�)�vQ���`cf�M�}���Q�/�d8�+)�/]���hfi�zox�Ϥ�c,ą�]L�`A��&���|��5i+m�_��o���א�qZ�������J�����>w�I6��ؐ
1t�=O�l���������ۀ��Q��3IJ#�ӽ��\k�b����rRϲF����fλviȌp��gt���I�.E���!^���"�zt
�����g�w��@G��v#6q�V>������Iߍ{^��Δ�<����h��yŠM!������(Q��E}("�z�����L��q�lJ��'"�v0"G���gm�+�pC���;�jTx��G�N���}l�Y��w��2�0�;��RF�����;f6�S�G|����ٗ
��^�� ?y�̈<&����r��y���e2�U$���U_���4�*�
,xH ')_��N-� dՀ^��vg�����!]���=66K���]���A��n|�9т�R��	=p�8'Ѳޫt��W��jp��u�d*g�Qh�M��*d��42�n����쓌���
-��ܿ4�>
�"OIȆujp��/�+���@�eJ$?.����u�n��J?P����z�͚΋�ss�o���T���ٞ���k�����ބH|���4Þ�h�,�#��ynL�q��A�`E�A䛵ܪDUשZ�8#Y�z��O9��+d�N}3:�R�p�|y�O��G[۶�����<�B^>:��dxБ3�����HW���S�<|�^���<�-F]�SϨm������"Co9�����]���g�'!C����X�����o��=�AQ&^A���8�ޥ��}�pN{��Vo�� r��@I�c!���br��䬛K�6�H�cb@�NS>�?cոx}}�уh�]Z�vGk����^�)lk6w���!�5��2Ic�99w�u�@rU+�g)�< � ����fGu$dH��_#�Մ[��OP	��`�g$���?�Na�r�ƿ	of_d�bVu �M�:�lK�aKbMy��V��0U$ ��f]�¢ϡ��p�@���6!�V�>/1 
O!;u����?�vV�A�P��']pz+th	��5o��B��l�P�ސ��58{�=醻[1��(}���!l�@����cY�3k�	Q*�KK?��1�d�&`�g���F8���)��?���KP1� {��MR2���bIz���/�"+�ُY�����^�M�[Fo�{�AQ6�(�oi���e��B?��o>I���*)��.H��aΑ{(�=$BP�8**
����޹�ɖ!ݯ5��@�9�>}���}��,�X�y#��.qz�̧�OE���jI^��}?���x�Jb�Q���@�Q��Ĥy����Luj��?����NG����\��r�$1E���"�O"4:�>���'�q���k��C��z*�l�2S�����>*Sǐ�i��-]o/��$NE3ػ��7Ф�+5��2l�x�jy��EF��4�;܂D~�vf�W���呺K�ٚ!P	���H�A��U}į��G0�K*=��}k���$�x��V�y�KN���=�)�����X���%�5���;f�c�o����J����¿��z�N�����k�g9H�!��R�/��KqU]�3b��w&��Z����Р���X��d˿���s��Qo8.h�9�o�֩��"�!�}����k�v5��1d|ωEW�W����E�	q�!����l�ŀ�=�_��u�%�":��dh�������B%������Ym��>�/I�̀n�ݔ���4i	���+0����D�'*@�����%���gL,m��8��
����d�����t�f����į�cüe��	U;�إۀǲ~A���v
Kjդ��ɕF�G�F7f�ҏ�	a9D&��W��͑��@�O��+.5N#-����n᡼#�gQι��;iR&����9+���*#00y[~7�����<�)^��k�ޮ������d	W#�Ҭ���*�>�\�n h5}����i��m�|���Aؠ?�F�G��� ;���8ݲn���-˥����,U�,��w�����dj9���aai�P�N�&��2MC�������,E�����NxlA��HH�>�5[[)pz��)����w��m���g�4���&���%����eŞ��g&-t��6���������"�P���Ba|�D�'7N*0Ա���/��}���"�:r�Zo����^�a�
�@�E.]���ہ�ޏ g�}��^�M�O�����˹k���8fi�ܲ�O�5kY
�э�/�Y��F?<;(�դs�!�J����'�/q�:c-�>�:[?i�6i˯v�8t>�'��gs���Dn� �&��s��ڐY�k�|	����5�I��9�ɶ.;��,Ňo�S:�5-�뗹8].�goO��,�����^�<�ey��ړ����~�]���eYh�t��n���hj���/_��ez�9!��s7�A3�μ��{\���4��g�7R�xU��6k��\��V _���,�4SP���`�yȒ�b�\T:�K�W<�nI�IHD�3Y~r����ca힋�}(����TV������t
���~�P�P}�u���oa�W�O�ϰ t�<|�����5%?�5������%���}�M�k=�P�����m�+2��������i"�^�./V�'���؛���o��;�_��4�H������f����:�1�["�k1��X�{�s]_
�e�ۧ;AL'm.�$LN�I�[Am.QBK,i���mwҬՐ}��9�����M^��ꓜ�(t���}l�3 D�A���� �i�Ub��j�����}������ĝ��-c ����p�N�D�<����3<Zj:~���sϏ��?���E6Ndڎf��N��x)OK��4����7�k�o,�f�ŇG��"�ӿ��$w��	u��0.���}�Ԁ�q�����F��'�N��@Eb:+���](�������+�h�o
Y��Y��9���is�h�5|������k��NtR���ᡫ���^p�ʖ�*g���r` Ï��l��Td�ڈ� �` ڳWI����9
�(e������_�%��β�i_�����l���ƙn)#���`���
�|�#�!Ig�5���N�e��ޘ��qM�N�p�=$F���_j��2o_�M�/p���y�SFi�wԈ���u�q�c�ј�A�p;ӀR�S2pl�+L%@�:��.f�l#�����鮀�( ��iC�-��}��B5S������1%�ʲ�[�t1�`}|��q�WI��Y-3n�oI�hڿG�m��$R�kʪF������>?;�w�����sx*���%�(�u'��I%���S�R_�B*����{��4O�%ݘFmo-K��?�&���?���\-��-j���;�)��q)2E
RPh$:���:�Az���>���M4]��#�3(!֛�a���L�ՔH�V/�lu��y��bn�1�l��sS��\|��ac�{����\��c��1�RΆSU�uS�_��8蓎��r�)�A~�.�{��<�tn�}8�M*v>�T���P��<D%��s���](�:��̍�W�궰'D��ʢ���v{��SGT�#��Sm�EC�p�2 ���|.�B�w�(��Բ�)Sa�툩1R�/j�kQ��NF5Q h-#.N���� ��UE�U/��Kc�A7N�Ys'�
Ǖ����>�A�?�C�J��(DpL}��uʭ�t�;C�=6f1ss���$r\���wZW���(裒C|!���zm�I��v�F��y�dK5a�tiC�� ��Y�ﻹ�	;�rj�#�2[Jf�a�#$�ȧC&z�����o%hొsq0�{��/T��'.���~D������J�A<��a���?}��{�������<쉂�Ee�`y�*��-�e[9�b/M���߼۩n
}\��a%��OD�借V-{Euh�.UI��
� �6�R�<9w������H8c�,f����ɡg�3âUS-'�ZhpD��N��b~��!|��'�UZ��b��NQ�*�Cs���ΰ&B�*�ks, ��%oo6����a��M�ڣ��r��qc'�lgCRT��K�Ñ�v�"��?��S�d��X
 0?=����%J�#�g��a�y���'�!4򌋏w�uK�#^w����?fVFl+�,��H�J�^��.;G\ۂ�~�n�%y��@�y+>K2��{�ZX��m��`:�[1����樦�V��S)��w�����t]?�G^l����~�NS��S��sM�a$G���F��푢�pF}`M���t�[�Nٱ��k�Ț?b���BK"_a���ڡ�����|�s#i`�&.no
�~�4� j��"]_.zI�]`}��|���2���a~�h]�z�A���c��W��8�	ׯ$��T�F&���L�� ��V(�q�Q��Ӡ�`�?�&���f	��(^_d/lXe$�~���#q��>�h-Rd�ޠ�Q�R��<��5A����NYc�Gx)���V�O@���A�w1T�Ǟ*����.������߱�i_?�-3T��PD_�NU�������V������AfL��H�v���Xib�5 ���h,fۣo3"��bzFz^Ѡm�`9�	�"��Zؖ:{-�o��������G��&�BU�TƱ��ܷ͠}Õ�������d:��/�*�\neW���eL^�ĭmh�Jq��/�s{D�Hiz��v*<A��_W%v �A���ϐ�B3�j&D���;V�y��7�A���)�?P���/��|NtX��6u����
6l#���(�:��g��qX���ͯ�T�]�5�d��ύAQ�\� �Z4,sm��=��Ab7��R��j%�1�J���/�1���mAX��z��k?���t�F%_�'6�W��8�"��w���O9���ޞ�e�v{�����au^*͢���&��f�K���?1ahs�����렠ka[v������GJ��������2["S�/S����ݫJ�[L�����d��T]�ȭ�WU�0j���0�f�Z�'�H�lnņ\�����V^/1y�U�r�� [�%K'A��C,<�伥4�ew�c�U�k��A�7q��Z��䯷���T�c�V�y�
��.�;�h��#�P�J��I�4�z�܁�� ����qQ}���0�t#!ݠ�t���H#�Hw��4�]�4Jw�4 � �����}��f�ٱֳ�z����l�[{p���lek�!�_8����ym���Bq���,�"��vr�M�Q�|�U���Od�h\ҧ��Ӣ�̳7�*5�;dP����:�v׹�|od�|n�ž�e$�~�"�1�qw���H��>��j�#��J�s�E'��~T%}H/���56�/�=��2�����wL�_'}墄��C�F�ۨ�I�@���[�w��q��Nb���[��麱s���H�z���p��/{��&��P�09��Nx?[���J�6�� )�$O��#K=�M�C3P�r/�n��:�ov7��cc�n��CD��u��v�0�^>)��gm�&Ŧ�=��0�/��u���4�7���^����#����!�6U�،"k�DC5�8�8����I�s����^ƀ��-ػ�7V�zfxt�}#S����r�����=���ů�DSz�D.ũB]T���Z|Ư����Q����^R*��ׯ������������(��ӎ�3���\ˠ�r��MK����2�N��Z��>>�c����߆���l��~3 ��p%֩k�o*�s89���&��A
�̆6&E��f�s8���F�J<gvҫ20���;|u�Ə�����k[�$��8[�u��'��:܎���З�Tpq�o)��}'B��u4�8**}�#��b�����u)�����a�bG��u�t��Ѱ���B�7��mS~>�B�+��g���@:��j��f��=���ɋ�'���>_N|b|�Q�f6�V�R���9T������g�8u�f��u�t��o����'O�j�s,��q����jvJ��%���O�{?4M���W�k������n��f�Ƞ��}:�o*�?�b&s�)��0)�/����� �}�o���H,�o�Mi��Gj*(C����u#�|���qGQ��rb��E��:;��۟�'�juY���)��h�������'eN?�gw1L��-LE���E�ZVð�%����A�8K��1����b!%S3��+Q�ݔ ��:�ηmd�7��"l-���ty4���������Js�B��Sx��abj���djQ,��F�Ij���f�$Ks��P��~K��_�`�F��>wI4�����x��|���Xϛ�@�]}Ru%p�e0STTo��pC[�5���׫B+~������eyK�vrC��n��B���L7�m�z�E�[)�WAx~rQ8�b ӿ���}pHb�ѽ����(~���o�#?s�s�_����X4��8�x�A�3SS'(��(`{(��y$D��o�\������]Д�t�#k���+�Le!�}����V=������J52�J�p���"Ou�w�~�S�W�q&'K�(�܂����j
{u:q��+ݪ���?��f�=R�tN�b&%��<;�������쩮䣇�/i�|�٠Y�`,BV�S�\��4/����@�J�o�7&vr`�m_�[Tebϣ�#㊜�����B��Zm(���p�)c���P�L1"����o���4��{�c8��N舀���&��h�4��T��������
]ϳ�{?�H_-50����">��.��&�U�%���� V�.�A1������F��.8 �W�f+�� !�u��j��^�R���eښ1�CB��zDf�}�F�7����}�_#�h����(�?���,��u�W�)���?Û�i��ȁ�%��B����{X�
Y�kʝ����M	�*_�I�g"'C�WWX�
%H5���i�D��PɳP��dfs=[�v#�Q���V Gn�u$�ß�@�I@V߁� �B��t�C�V@�n��xN4�j�}�w��o�;�K� 쌖����L�uqr�^6}�sqX���u�C�8s⿴������Ž���d��N��}�V�v/0��]Q��!fX�8TB��y5	]��ytl]m���L$˳��_���v7}��A1\�MX��Np�SNNƹ]&�>Q�|�@i����L�cZ�qSTY4)�Q4��3|�5��ϛ���}�'����r�l��o��\���ڻ�ϡ�	젳WFS~�\a�Ls�#�q�ab.��DcVAe<�q��-��%I���,Y�z(��m΍<�wC��~v�˃ H���|�a�b��,�����|�D���"��=	g����_1�z�����ag�k�X�cI�q�w�����w���e2Ɵ��CP�.Pܗ���R:�:�] ػ��9g��lh�^���uݞ�����xξ�Yld*��5�$Y���%Q�p�����G����־� �%0Yy����P���_��#��d7��!e�["��<6/�����Q��A���~Z<��V�2,&��d���!�����}E���'���s̢EN���Ƥ���t �D\؈�n�8y���"d���>[�l��2TJ����T�c7����_��=�d���Ol����z\t�g�e�]�R�� F�E�{E����GZ�w�����*�%�qˌ��9�T}����9^������aR6᫠�Px�3|ZW�]¼�d��6���lзtx����[]��2�G��q���w�
���}�8��8M�	�:��Cs(Z�����J���������\�=͟�m��.�$(���|9�Y�8��yv"��$m��H�w�Tn��E~y�~�5w��~cGC�<.[k>�ٻhh��~D�h��'����T���K7�Wj3]~]��9���hr�W�D�kc�=|K#x:��S��N����,�Ԣ)����Z]��T�6�b�XҮz~�S��z�_�z0�P<�"ˍu���t��q�+T��HϾX�77+�ǿ����M�8��s��p���_]�=x����!j_��rr��/�fq�s�"MՋ8��:�A� 1���#��jƼBA.aj>���p�[;?�����B�y��
Yc|o�oWv��JH�	�����p@�*�����?�}p��?F�N��?U	 ģ
���13�w(�7�\�|�{I\}o��s�a��{?��9ϲTW�
:`{�d����b[�f�"�NN�{2���t�'5������;8�^�����iT�8�O����b����;����Yׯ;�9%�Xy�̫�GY�wa�����O�Tg�q������X�t����{�!X3�N����yyעZ^�Q���9H��R�ٍof64�
�&�T�ä�}N�q.���o�t��E�P��j˓a����n��6]:����yN|�f5�z���[u��[*�F�c��"����Otǳ�g�8��gOi݀W|���
�������:�<���&4����X��EV��!c��������R-�V��U����������e���1g.q����N�S;�uRW�nu����E�Tz�R�+�7Xܴ�����'���L�(xE�n��&���3�C/inGJ�A�����(��P�RGGez�~�60^ͭ��Q�[t.ѭ�b����Y�!�8B��r����	h:*���q݅�v��*�*Ǐ�)���j|��Fyu�9𯚼XDt<��ф�+���}�%��񚚍"��Η���;i����a"�i��O���ʹ�w���*��H�1~�ڬ�[Q���,�`l`s��"P<"ݲ�'�Uϲ�����FPβ�d��[���Λ1��Ie��^�O��o���]��/m�Rn� C� �����i��d�&���K��`,!��۝~ߕ���_x�7�D�s��Z�\�>�?��mj6]���贍|���ﺁ�̣�`����^p��{��q��s�IX�c�����!�ѿ#�˵�n��L���m�l�������j�ύ�K��� }���?w�f�(���� U�������F��IՇo;>z�/�jG
��eW�"�(�ē�+Ƿq�1�+,��-��{�v	��Ff��C����a��U�p��P���O3�2V	]���"��F�~Ss��?�x�?����䒛;�6��.L��ݡ1�f�*���*膾���oL}X�28PK�s���0?o�+�`�������d�K��XY������Cz!��8�������A<�nX���@=����*�kab�N=FW���3| Ō}�h�
]Y���>ɸ_?���S������b����V������Y��&x�˼���ۭ��u��ȏ �������Q��Ǭ�a�W��Bg7���s!�3��I�W�c�kc�8�+�Te<h�R�BcU��yd�Rfc}�c�$T�DK�4���l0i��g$�<]ot�G��*�.O}�x~�z5zo9D`�Ġ`�Y�5z���Vt��YԡÄn��Ir�M��1���t�����tZܮ�*���P
�������J�h����Uj���h�!��CL{�:^�C����gl���}��rSr9��N/N�i^HWc�RU�`�8T���龸��
PY���|T.d&7�a��.�΃oIÎ�3 �X4Pm�����>@�o7w�������$����,��.k?��`�Cl��AX�{�3�/l��ؤ��H��0���d-��xy��K����X<B/wް��7+ϧ!�sx/l�Y�L�����P���X'2���'���9�����JI��p�8��˻J��+D�pJ��A��Y=K2p�(��꠬�HX�I�#�[q��l�cܓ0@�?(D��E�П�����A��\Ā絥�����o���8�ź<߾O��c��}'���s�E��~V\�aɮ ��pd��7B���0E�P��O�;e!���'r@|�~����w�yQŏ�N��v4����I*h0>�4�
K?$�ȋ�Ր�eZ{�?$�;��9n2�(vDx�>����䭑f�s��t�`�Q�:Fq(������������d(���������	�cH��W����3)�X8_�7T�ܧ�,AIP� �:���j?a��� ���
`����S��I��"���)(����xe4��|����D$L�n��wn�Y%�����-|�i��\Ďވ�&�P<��`�[d~]{'�گ��1Y�"HY4xm��N�/h%ǁ�o/��.Y�㓲��,��L��Y���3G����Z�Z�2~0Alv��u�9�vlņ����`G8�G���zI6C�b�����{�K�?��Q�[qb��mz+�Ĭ)��?��aq/<�ä���X���I� �{g�h��z��Y�wD���V�w�g@��P})+�l�|a�l����� S��@p����uL�� �������"�뺁 �6��7�jN�K^c뀂W�f�Y��%Zl�2��R��jk��r����<��.I���*�-�Z�@y�d���I(�n{L�|d�8g%�[L����C܁�Ip�/T%Z���NM��2N8�K,�h<�W%��|u���I����â�E��;�/�,.�&�
L���S����t��.���@99q���̡��9�nIgN�Ӷ\�K�'h���kT:)�����#z���������?�g(����et���e[��O+�q����|�.d$�52A7�C�5�z�/�n10�����`���v[2�u�Gm�?W�uu\��E��"�+5��ÜBI�rK��~4���H*�)���J�W)E_نT��
�$�D��$�KF1���������m�))�xq 0~����ĭ���oC���z�* �>��(#i��i��,�~��.���p+��N��#���b2]�OL?�����ʍ�2����G�G_�o��]����mkB������m�%�4"�T[����u}-���YuR������9��
)഍}��[N�2�Mƀ�ˡ��~K�7lN|������7)Rh���Z��d�Ϟ�69cX��'+�)::8���'��y�We��*�������핀�j�Yν@�jYt5����Ǐ{*hG�f��EN:�Sn��ޗOQ}����;��;>1�#O[Ky�hR�G	�]�}T��d��v*�7G�y��z�BC�s�3!f�-�{)�xҏ�tL�@-��Q���bO�}n���.���~u��8������eaw�٧o�Y˾z�2\((����u���Q:*�4�4�y�ʴ�k@�ǲ��`:��q��R,�����I�n��ص������^�1��έ^�bd�
�I�2�~ms��Q�JYN!�Pe�ʋ��A?/>�;tT��S(?���t	5�����9	A�i⎫�(��Z��W�㠒�ā�Y&f��A�`�Ш�LM��P>/�j���qU�m�� �7E=ڭ�>�6C���i��2��=j՜�+�"d��vb�-�B�
i7�=���1�l@s�o>T�y*"e��Sr��!�wjf$%����O��Zu�#ֿu.G�Z�WYC|�|��%��C�����U
&�w���*��&Сe��tn��}�E��	��R:�-ɗ	*�yK���������'� �/Ǜr����L���#R
O�����e�˝��g�r����ٓ�T�W��'˕2����F�B3y#�ux&�M5(6q2��r����*���F�˂̡dn�d��3ˬ�6�� �����I�W�N�����0���M�h���5qr�M�:J�'���瓙�P�)�4{���=l�t1���&���Ԩ�H/�����/�]�,�������a5Gp�@�����j��zꢲf���G���� H�|H���ӛ�	�~2��5�ɺb�wn)��(��
#�륈�S.�6�>^��n���(u������kt+}��M���,>
����,(�{9��7�K�YW>����ײ�Z���):�)�W��q�5�L{�`Gw|F�X�E�<��yY���=�L"1����aR�m����a2J'�����Su�f�/a�=�c�-�q���{�� +7�_��.B5�7W��@]���G��ǡ@�O �ON�Ĥ����'����I�����9�V����C�Q�-�-� �������0�v
�Sֻ�q�����˪����J	��c�f�!�J�-N��`����v��I������&�1�'���
�M���{�{��]�o{Ȑ2� 
��N��E�Y��t$��x�N��<�A����M���/�ػ�L��>�ɑ!J�n:�--e�rm�3�O����C��y=H ���jdR�ϻM�9_���KMf�k��i���I3�V�p���r��p��D�ߡX�\Q4���kOYY�r࿝�bZ��F�lU�i�8����9;��.BU��[�$ w�42W�٪�&�+�s�J��#�X�������f�/��* �UC����Z,U�5>�1�w�n0^�O����[:*=M�5\h"m��J�e��++%��t���t1џ��d�\S�ȅ�
4�ԛ�`5Nb�G��LP5bw�������{	Ǜ Y�+���q��W>�ш�Ox��t���\�d&�.�ۦF�iab�dy.$��B&m#�*��q�b���3�2 Ќ��G7��AObȝ#(-X�3��hGt�UU=�n�r�ƀ�����_ޠ�ℨV>���v�ة�[J��)� �-�_˰7�q���F���L�2�r8��jd����3S#���	6�J)тC���?~����2���ڱ���W�ŕ�ߟ- �M�vQ�-�$�k"���dc���V�ˍP�q\7���a4g���ptk�8_KX��6_[�8e(1�/,ԙs�p�BB'�_��g��ǡ� ��c-��f	E�A�� �@q�t�&��6*f���vq�鏌�����lن���У3����{�A���
,�aG7�:�2�/|������Z��ZR9��C͋�����êO8�X�K<A���Fp������,�����5P��V+'���(O&�bNhP�d�6�@�o� �y6o�-��iD��"��{�-E��\r ���ع�FHe���O>|�טG2���s�D>_�u\�_��A�,^��n��ĵ!ff=���b����;ۮ� ��ۯ���P��Cž�WӮ�Jt�	�R[��e2�]�_����h�WU��6+B6}�<S):�m���J�2�?�>��A�ؙMp巣��D�)f��������&I�ר5}�h}Xnu����G��ߣ@.�(7x	�4���'��p�:t�_��q݀�4D�`ڕ�(����RW;d�̌�yX���hX�ZUP4����S��)ftY�4W�Q:��ר��z��"O٢��foo�����y̤c��
CW. �����!_
�+��j&����MΠo!ؖ%��Í;xE;�&3�>�Q�e�II���>Wi�Y\Q?��μcukS��es�wS���z-6��A�g/9�d��N8zd�~hٽ�xx��@���@�(�/��P* ���\���QWWd�(D���jХo���ػ��ms;�����A�����/�98t/�b3��Sy��E��jo� 05�AJ��l~���okuH������p*o�سﲜCc�1˹����ǿ#W3Ks	�"׳0ww�j9���&r�B���hݚ�D����Ԓ��C��"i{m���ˈsYlW��d�N4_�9��KqX,�x�49"B5����N_ʹE}�c�b� ~�#K��C�RU��w��
W!�x��p%=�9B<�a~��r�v0Z��29ۀ��ER����F����
�؃��4,���ߺ����kKx �ŧ�$H-@0ݎ��܈����=�����nFO�A���d���7\?j��y�
��8�̆��`�H��������M�@���m 0jd�@��	���� �����ueE|���ĝ@��!*C�H���'C���q�a󱽃l�V ��he�j�E��Y�*Gc)�.#�?X�O ����"J�R#�߶(�K���FT�/҉pOS�t#)K�T�����l�I'�WY7D��x�iC��M���>]!���P���z�1g��4y��!u2::࿍��<ko���`��l4��
I��d1�0Y�c�S��(�\�J���W@�@
3� ��'��^�k�PßX���X( 74����f��N'�ۍ5����L����:\LN�j��X�rYQ1>�^MJ��~�F/�֏P�L��kj��C2C��EA��m^5��q~���!����a����Z���ӕ��斥<SD-�f?�r�nZ�7��94]�B\:�2R��,k >3�!$T���@KX��3,���R��p�����0�m�:��fK��c�Y�����B��0�^��x#�!�!V�_��M7�|eQ}n�w;|5���kr�\�|�x��JAE�C�k	�C�:9d��Ԟ����I��x0�B �,���vÆ�sX?�Y�Y�v���O�f]����:=/l�x��:������;��V8E�S]�j6�W���y�̈�F,O���+�J���B��F����C������p�E�B]��$⢎K-�Bw�*j���I�YUJxK�����K�x�5����;���|�ߤ�M���ݜm?I��l��KԝCp�X��l���L�*@�����e�楎*�l���QPsl���_��;G2�'6C!�w�|i��շ�x؃��%6o~��MS|��m;�J(�D�H�!���B�m���W+�\�Tf��Amw��K�2��|�������"e�,VB���i=T�G�%�J	4b$���2���@�u�)�_�4��9t$�x��K�C�ZJ��+b��?w�pb����wI<-�*�	Ke�#;�U�]֡��	(0?2�a�i;W<j:�X���b�+�t���e(���i�GC`>�m�$z��<V�su���ܬ|�w�L �/|�>�6�&h�8:Ė��qP΃������1*���(�0cx��K$%���%s�N,��xHR0K���z��X@c%��O��LB:�%���(����f�>����Dbe-S��(y�?TN��!?� H��_��r�}$�Lg��B7��A�-�F�uW
���Ǩq�@;
̶�� G��j���W�&4s)r!�SiL��	a�M�U�k6C!�9�9�O�/#�ҫ1�Rś�{b_t����y�ʡ����C {�;?YTZ��Kc��!�	�/&�5�x��+���6�k' ��{���*B�Cr�ρw ����:C@4O����iI���yȎ�Js�"�c#�Ɏ��
��r˻����2�����M��_}�j�cP,�/�M�J�IH+�G\�\՗С�YF�R8_V@t���uE�O��eD<6��'x]+�d��,�&Yp�x+P�fN�̡��}�{�{����&$��,>�����ǋ(.C=J��|y�c�y�?�(��eu� W���4͑��	�<	9�����1i.����������_7t����uYZ�׋thG�}�&ȝ� i�RO�y,ܜ�����~��E��y�F�/,���K\�.�������Lڀ��A?VJ�W,P��ሴ���� Pk�T��uH�(&`���2h�cCH����w���(��N$�	F�������H"�n����2k�|=��u��j	�����fT^r����w_����%`�������P�WL�@m9f1��ͪ�G���m�u+��EE7�,�T0O�]�Z�v�`���i�~�|C )0b��!��0|�" �o�ʡN�R�,��aM�p:\�O�������p��\���$��q���1:�m3=_C��Vg�����  /9�'z=� �	�=_@
�0 $�]_�,*�6��eQX�K�^I��������dYol�:]�9��������8D��,~�G���3��S�ϊZ��q@|�0Q� ���}t���Q�����/m���r�uv%B�ri�>nB��� D�ģ�6ߢ�@N�o�s�f��MK]ث�#?��7*ʱ��y<���I�0��0��·�;�㆐�|� �����,��^@UC3U��4gn��K`�*��Y( ������y��x#1HtAUbAԔ�&�q�{m�8(<�{sH���5����a�ׯG	�D�e IUy�<�NP�q_�^���zZ
j��/�UV�[�٘L^,�윓)���3S�8>�Q���T|�0tEw�V>*nj
���iL�N}�2�ɿI�gL�����E4��	ȩ%,~�3(Z�bR��/��B;���X����\
c�͍�#��H/��?&��B���;�4.ĺא�`�,�s�!h���@���W�o����׾�c��Bѧ��F��C��Ƌ���ۼ�$K+uAo�}��įtA�#6;<!?������	���o�!���$�t�B�)w�'6��z��ɏ��R2`�UM�b,A0%�@������nҋ��>��Ht�r�NwԀh06q�:�r"�Y���)P��Yqk�\1����>��=�X����.D�����\v _��кɑݻ�]��
+�#.�pǛ�51S�u�S娴P"9%1��m����P'��&i� vv�Y�`C�R$ 'W.l,C���w,��hu�g�>��4RgpS��bu=�"�
�8[X��c�x+��ڸ��*Ǥ%fl�vK�* ��r_߉E�c�2����=��h���
��kni�'Y�'6�|/�&\x�����+��];i��}�|M䷧�aȑ�t�n\�=3��CX�.��� up��(<��:�@g���IigjP�ͳ�������ʟ`, ��	ts���8&��w.����K�a	ͬ����g��YGG�O$�p68����r��k���C�*=59��;��sL�c_c��e	��x8?/�����:[@��^�a�$ht��HS�cN�o�����#6�&�h'�\���?F�c#7a���}���n �{C��+���^�(�r�X ���h콻!��!���B6v󓞟��<svAy.���-Klդ���!��β�����O���p�{6{D>͗Υm��3�|���YAq��Ȣ�P�uD��i�Ħ^B�A��\��- �)�|�'Zl���uL����@���p�t8B�/n#�b��x�(M��r�YOd[��KS#��1���۳�i��ށ�-r,$%hw��Ԥ7!����F��Ua��G��~��S����!kEK-��!��B�-! ͆�X��RM�گT��l�; �h�`��ի��k�n��K�榧q�v*�ʰ��)S��W�W¥,�����ީ�|aw� q�sٰ��t� R<�e�V���yy�s��|P���5{
H?�����%V*�1-�U�JJi[��*M到�x��c�Θ�ʕ������|�x�'�S��o	�7���YM��s����kf��j� �H�]l�3��C��+�1�����j����������G-��}	L]��!���J�2��/"�6�KE|1W��ũ�G��"�-����%�3$V�G�.���-y��D	�y���CѦ7���xd4k �ۈ7t��w��
��+�G��(G-fi�/�f���@���H��G
� R2��h5��9 ��6P7P��Ѐo����m'~���W$$)�u��
�D�0vU�ý�9�yj�g�r�wO� )Eac�?�>�Xߑ��shf���
�K��J�u� �pM~f���j�'ɫB=rX�4�s"��u�|K�e�����k�S}�F$�+�����aE'f%e��y�'�S����4^<�\����t�|=��p�G�=q�"=���S�?զr"�E�IC�dq����9@�M�mUkO�ԹM뺕�B{���H�:�L��n�Ef���e�����_�5)	�F�d�?��C�gD,]��Ƕ6�tVw���[���6��������H�$�oX�r�qI`���ç.e�Ʋ挍-�w_9���;�^M�Lifa�/�i�#nRH�-����ѓ��A�[���J�^kC$�]�
=�7YWLUӘ�a��oe�b�\KE�h�l
��jV7��(gV~"n��Rn��W�H�ֶE
چ_2+)���Ij/��K���t���Y�\����Sg=���|�.���+�է.ٚZ�7k�0A/� -4�i�mV2,":_�������Ɗ��kf|�*qw1�y�:�r,��v��ݔ\��}�P����g)Hj�8y�6^�e�-f�9:��P�vR:����@����hQ �_ډ���4�Ц���Aj&ס?E�e�j"U�;џ����e^�`2��8�*b�Z˱�$V
���K[�C���!��>�ޤ �+7ܿ�Y!=�P1�:��{c`���ݭ�]}��[B5��H�v��ԇ�t_�D��@�lQJn��ŭ
��R�Z�����W�H���-���OVU�֡����BPU`d�|z����8(���0p!/��ͫ%��a�T��af�Ӹ���aW�����x
���ul	��l��&��z�7ӏ��*����k��%!Dk��|��b�v<o5��M���e%���}��|�&Q���>6��ئ���@zM���\�x�ݞ�9��(��,�ߦ��]e� wц^�D?o��c�v�Ґ��h�k"P/�7�v����������X��)�D��7��tm����U�˩�|Ǒg£�%V��T�}LT�xB Am��G�-�s�
t�:a!�$��N�Q5����c�$�c�a��'�3vx�_���͹e_�B&a���>�<߶ P;52+iL�ׅ�N�:�;�J�������%;��������ZNn�c=���3���i(�� ����� �E�{ns�K׿�Y(g=��3�|�X��;tK�ǡǪ��<ou1��ܟO"���][������l���G*X|��pZl����]���z��Xq�N�ٗ��%U�?ۨ��W(��ܨK�k�`~3��6�czI�f�?5�^�튮:�4�v��9`�h������{����C�d�g��+-�yB�\�N�`D-.�>�Q���D����TKKc�� d��H�Q��n��3�Tc��R�r��}���u��h��ݗ$�P���V���?�ڝ��w��ɭ�Y\��h����V}���������P��"�
<;pq�4�<�#s�G�~�U;xMqҁ����]޵X'��{�*�����5�f<&��ӳ�.�{D�ߕ-?��@�9���n�$<�<�4!(I$؄��XSS���<�	R��R��B����rX{×���9H��츊	�������{/��Gh�@M�T�cN�X|�@aߴ�����	��Z�{��L�?�0�O9�+{ɟ�Oph�)p	���h_�bj���2ϜȠyab���c�)S�L����+�SK��V�Ч����;������)��%�z���#��5_D�l{TWk�g�G�罉������e�.u�i)qKQ=h��3�.F�@c�Y�[t�O~J�R=���4\�=�~z�J�x���� �Ϊ!����֔�e+3o�˃�`��͍Q:��\�9�^��2 ҂j�vZ,h�(S�� :La**�>0�8�#�D�nn7SD���Ֆhq? ��,�&��,�����?A�W��,��K�i���km��n(�)�L��ğo�68�KP?��+�Lݨ#t�*�yv�d�3��d�oʫ��5�]���V|���(gbJ�!b����?�d�$��b�.�^�$�;��Moj���C���퓝 �pLr�r��%�3�6�L��� \��,�n5��h����]���>6�d#��%�>�3��+��W�;��O|j�R}�4��[.8�bO(rӺj����S[N��t��O�M*rs�ʖ'"��Y��[���%WSD(��uocqg�L��THP��ia$3���ֱ݃BI�n��H!^�㮓$HI����iP�$��sBx��{1����{ϛ������}��gR���k���7����ti����N�X�� v����3��@��������E$��e����Ԇ#zY��=
�8܏d���[
�?�D��mY&��dD��4��ob�ί����rHx��aC~ӯ|Sw�eq1�~Yg>��uMy��׾�,��lI/�6f�G���I�Gdw�����z^����w��mM�r��T74���u>�}�o��	���X����Z�9�SǪq���V  � �cj���;dqݕ�g����q�hA�K�`�\����i �Q�V�;�������04d�X]/��I9�x�ZK�w�	����&��@�k��$�>8���P���;�{��b���8����0��+B�.�`�<_�I��}�{�9O���7Y³�/�8A��u��)�p����2[�|ۛ�A�Vɒ)z�SL�<�;�� N�G(1rp`��8����Z_�jw��*Y4i'���Y3j:��/��$�-�#*�� ��M#��޿0��7��[����)��W)O�h2�|n~0�|��Q������R�^r1�~79�,g��O	�ykVL'��c�ύ%#A�	z0vF�Iix�392�κ��W�;M�d9���4fHX�x����Ɲ���L��9�q���F���v$CSO�+�����;3K�6X^O�v�ӷ���E�b��א��8�աc�OOlVϭI�,�	'C�5��߇J��2(���e�͞��:_�r��l؇�I�Qg��,�3 ]J=���
��UƏ<��xټ�f�IJ����R�d7��9ږ���h{��δ$�SdK��<�*�"�S"�A\�e򛂖/�3^ h��+:�6��#u�㾱�y��m#��V��Ұs��?mlsv �t>sQ�՚F�ޗX�/7�;�P�<>�w�	��e�&��H%{/������(��B�__X:��ಌ��0��xȕ$�cI����bJ�z����Ç3�k ?}�[�@΢P���fe�?�*�@���R�Gw�.e��RE@�(��f��9�S̻W1���}y�Y
Q�xp�:���:ڌ�_�m�'��_^�i����Ѫ!��n�[6��?�
��H�j4��5�?�� |����7,}�ʡ�ћ���E�or?<2�����SQ�=$	���.�cT{�{�~�X@Z��Q�)���E�-dO���X%��x�W��<���n0p�$7�c(?��c�����}`�M�_^���Y{ �ɲ�V����֔��V�c�[����%�]cM���7��U\^&rZ�><��X�$��V6~�k�m�{���I:L@f������V���	JC[[x��B9��7-�q)+����g��;�PƊ� l{3��^�yo���m�!��8�Ɵ|v<�4 ĭ(���*Wߑ�dnT��Lf���5��++.�����oR��:�þʢn���0l��[���͏�/V���w���6gx�m�	&��y�[����k���>�g��a�������D�1Ϊ�0�?�j��n�Qf�w3�ʮ��!2%Xէ$��2 N�$X,�����[G܍�W粆��#��o��J�ܶ��Fv�R6UE%�3��<����0e����m�y�U�Y���P���@�{�!{�z:N�@F�9g�H=����;�]���(<�����N�Ge4bQ�I�����5�/�H�ۘ��A��Q�h��@+�T��v��wE��f�5��-S(�`��r0����8�$J�%��!�*���S\M�5:�{pww�w��\�݂$�;�݃Kp�!��������?�V�S�JR3�{�����9ӃG=|� ��q� :�NǛ����Fc0�f��>$9#J_䪼� ����9�jғo�M[H[�L���>ETs��Q�~> l,-���/d` ����"�oкՂ�,4���#�>9~� �Ȩ��mк�6�ҶF{[��K[�/��G���ɭ��&+�N�E��yL#F��r���R݉'4��&�j���}iz���sił���3�G�. vѯ�?!�����Bf���Z��{W�����z���:Y�t���p7A����z�1�8�&ǩ��t{c
�U��g
���.16�0��Ve�����4wH ��#O~��u���F�k��ل?����p�g���1�՜�_$!_�?`���6���[-x��d�z�ST(��%^U�9�&�Lw��Q��1�����&�:*=����������WO��exPv�l��ޗ�CT���xs�op7򴞝�U����M�x�~�z1�����JXFދb�'����Z$�t�=�`]�}RwG/�;��>o-���)ԠyY{�]�LY���ވ�R=\�0ZKV�{mkί�o'�c$6"|YJG�V��[��Nb�L��B�sV�����˿5[7�E_�G�`B؟io�(���~n�;Ǥ� Y�'���~�Wѩ��֒u�R�|��i띔�D(h��C3��/O"D�A��ƀ�5�Q�PzS)�`��	�<��\!�K�p���^�m� �Sv��ń�^g�N:#F
�jy��;W�%�q���X8�&#G�@x�F֖ݟ�O�Xx�V~Ub$�h�z-I"�$?{}�x4qLˎY�IC���̪A�h��<���ѝ���	��q������i��2`B�h�1&ˎ�笖?u�*�E��!*�Bd���J�W%��ʬ���=����lR_��ڴd)��~{��!��u} ����S�ma7Tj�́<�F��d��l���IOJ̄����;�6�:��Q��,��S��Uo��<�6�~�	L�{J������UI�g˷�qId��_п�¼'��`)�����!�u�K5V<i�����m�!n�������J�ۛ:�(�.=_�G*8��E����rj<Z�5���6xr��iNѠt�SҪ�����&��~֪���{�F�P���Ni�Ռ�^�G���Y�ӪD��r�z!� ����D$8I��Q��mKY�N�-�B��ā�V��\$�<9�̫_��C-T�5�'�BYao�޻�͸}^��x�{Pw}�*}�t�T���N�L���Z�����E���*m�7�����ᤵN�)w&����{�}��;fU����6�%\��9\6�Dt���b����j-�.:�2�V��P�F������<g����)�A�!\����ϔN�\���`ժ뢥���4:�9��G����/JbD�cbH�&P��W���D	Ŗ���JJ�\�F�F�I��-Z����J��I�k f;�Mo��>!y�`���TLf�>'�94h�lP������E;��gT�"yf���J�z�/����)�N�du�7�����;�YFX~��R�҈���4&��nq��T!3smv&zf�����:ܾ>�lJ��JEc���<s\���<'�����H���xc�
s
�Tm��$X�0D��;���&�Vs��?��$%�lV:a&����>sb=��=z�D#�Yj:�d+�S�o�~���3��;�,C�"b
�]|x��e蒗���%�� EƂY���	>Y���a�e�Ņd�6����7�g�^#_�����t��m��[M�Q=���A��	zOe���4�V_T���3{�i��4wC��Z�"э@`_
�Y0�tur��?Y�<Y�֖g�L����zy9I$��/��F�9�����d����%lxNo�=����W�T�M�ǎ���h�1��@ҨR_��f	�61����y���=-�?�&��rV�h��*�K�:�,�^?|M2�mM�� �V9v��ѫ�*`Dr�������yz��Y.�Y�W��x�&��9�w�0K�ռ2\w�nH4q�Y��
$'����(Z�V�"QG��2Z�5Ԕ��O4Hw�x^��LZ��I\JRz$VR��:�����&���������]�����qfT�(��$H�Uڤ!rн7�A�X�Q�۷+�����Rj�đ��>��H~Z��e�`��<`X 9%�~��? ɾg*���S��H�*w]J�ND���I����'�m�)��A9ip��JL�h�Ĉ�����%>�y@@:�4/���r3@	���\+D�-�D[y��溉;���Ut�9Żp0ɵ��R�A�S��ʠY�����]k�ߍ���w��.�,Wä��g�ǚ{~=����Tۃ���h՜�>L1��.��B�l`$��5D~L��F �w��)]z�3/Q�����\��*
$2�n�*q5(�4S���|�2�Q���SX<���
@g�OU_������9�����G1o�wp�u�&iC}�ar�b���L�wT�1�Ñ���t��ް��c%O�~)���x�>����s�F%�*�uĹ�	��(���=��}I�MFy��Jͬ�A*�,W?�����-]��$��'�$�l���k �e]J�1�rVl��w ���a&f���ǃQ��d+Wĉ[�V�ɽ��:j_�������}���x�"���ϒa��F�48�Л�"Lv�6ō(!��������}-<��,�×������3&l
�j����OY��0��o枾�iYSY���hm����uѦ��G|�1�+�1�A��y���Gg.���,��N��=c�S4PP�1�3I�����ͥ蒡�]�r;� ��z̲�4�uF{�~Z*܀b�np�"P<'���'��R����e��	P��O8������W˃N뜺����ä���Q���_��m�7�#�lf|�&v	I�%����Z����)��N�!��sn�D�rS����Z,��"��:?�`j bh�k}RL��>��b�&������mj��sy���9�z,�"+�7���12,�K��-@�ϤM��Ҭ�
�bx�%�W� ��P.��4��=�؏��@I���Ь�x(-��眄[6��F2+����Q8����YaAlC�\�L\"�=/�w9���Ttdz�ɉN� ���Ҥ��4.{1J���'w=_���5E���Nw<!��f����G�k�j!���2ǒ
�Ӹ4Z�_(�]N��
 G��+QN���y�X�O�!�\�2V#5N&_�іo�0 |�NEl��Y��4�$��!�*��
�b	3�����P��G�v��_�!��͵tA���/�/�y���k^��:
%�T�J��.�h�z��Xڄ�#\�U�7�i�ʵ����J ��m@���U�e	���n�I��;���z�}*��s$�º�La)��� ���|ǩ�#@z:x��}�ϸcZ��LB�Z��iZ��2D̉�^L
hOd���b$�
����HU#����d�tW�.�4���ezسY���I:����S���ضke�(��a/���1oj�]XV��g-K�_ِ|���D*�Ts� G��f���Ӭ����_��'�֫#O�za���.�h�|)�0Qr�g�K��Yx�E�ӖVd;Y�s`�aRhA����AZ�c;ЮV�#eD�o�J�+�|zʨ��Ө����*�3*N����L��=���Բf�aY��نɋ����Z趣,�ɥ��OMȁZd��m���c����tBׯ�F��p����Y�q���z�(wV�O^���+���Xޣ0˖=��z��g���6>J֮`9��E�qU  M�E
?�I�2��yO�T���m���(� ��r`gk)�Y�H�j���ȳlB��^`q�y_��ih�-WCa�A�	�z�qav�*���qj��v�DS��Ng�h$�� F_��^��6���r1tvtY�	P�3�	�z8�{�
�ś�c�q���ì�(�\�=T\A��t��O�L��?�d���?R[�3@Ub��)��R<�S0�(����%�g���Y���IC*i�lד�Z�V�Q����5I͌U>}��9/4�#�l�c]jl�{��%34�P^�E��u�����cY�V���a%�ƃ?��8��'�RF�;Яi�^/º�m�zg]�Ty.h�sb#�J�Ԝ�w��d5�>��uka�O�I\�崂���ia�4]kζ�'t�%��A�r=���(mX�	�ș�o�0��7&��(սb[�� 8���0Å�o���|2��8w��=��)kD��I�ŋ�d�����I#+��ݽ��e�����k	�͏�@ar6U�a��x�ìv����iC�� _.;�9(n��Y�ʧp]��Οk�����6kPh�"���V���:/Z��i�km�G!P3XX�C+�{�Ї`ghh~�d9�
a��%�q���?NR%W���1;8���%��A�����W��������x�e�@�C(��k�a�+��+����d|F�f�LO����Pg7}���-��èF/�FF�_Ү����nis�9QY�f��M|��� ���Za��G{����4����y&C�kmM��4�gF�iZ̮�k�V�Ƌ��7��X�4�������	J#¿C�������1����:�Y�<��P�7��O9���׺I�9(C�0���vF��
��$�}�8y.�����3?3��٠,�ph�Y=-IrԳ�5Z2\�#���6����>�����{��#Ɏ_ln�@�R����h3�?���_��[l}�X$9�������o��=מJ(˔7^2�>m��/��ԿV"I|gv~/@z�? ��ME�b���h�"t��P<���`y����ꃊ�w���e��R.���ŷdmkd��  �&���.�	'
2�b���L�{ꌧ�Y���L�7�(�ZpX��%����p�������f!����a�����O�/�����8�h�ߘ�Ja�|�ʗʷ��s�t�f�܅j^X�)y������NHr�<h2�!�w�+b(LDG�%�{Y͔[��~�p�\�2_�:%�E��r�S��lQ7*zC�B�����&�^��G����q����0�Fz��7�F)w��0l�GY`���z�R�@_�M�0�S;�����5Kȣ:�òtK��;�h<0�Y�S,�U ��(�x��P�&W����>r�mVE�ᨖe��f�;_���Y�.1�����R1A���l���G���|�as���[���h|�(�ը��܇�\׎��s�sB�9�]�\bS�l0pWf{�}��"� dF{�G�]\���~�N��#c�����Q���e��*��z��w���D5uE��f]=�W���6�9Y{�jo@C�8����������)з�:jg΀U�;��٫�î�
���ӈ=F����$.� �Eq��[�������ˬ=��0<��O�&��-�׳��7��w�z<XI�������:�@�Cݠ\KO����:���b�g����QO��c�8=@1�Š�.�H�[["ӧ\�����Xq]\&��w��Zw��7U&�����^0�xK0�'<�c�g��0*T��,�9��ݛ�P�4Σ��"玺���(�"�'�f/0Ѽ��M�B��p4��<���iR�����
�a���ﰝ$%�Q��.4���*�3�H��/?�ԄI���5�y
<��!�֕�;F�4���D�,A��FK'B'��S-�������>�ǁ��韗�T+����t)=V�S(G]	ͮ��+���4p��֐nB�X������n}ģ�5�J�Y���$E�������}�4����D�t�Mo̪5.��o�	l+/m4�)�����*�o����Y��P�'��$dJ�M��	�e�jN�x9ܝ=�|�QB��zQa�˂LL������c1��O�����`H�-|Ș:���p5�������}(���V��<o���D��@�n�|l�ykRв�bz��[
��'ʹi�=I^I��HV��J�ne�9y'r4�ލT�D�D�h���a<p�[Zz��Me��Q����]��{�O:��NφEX��ʺ��Yǂ����Ig���N�T�'��?V��������=��0A�;I��!U�{���/�^�d���2��r��	[���<���G�U@�i�A_;s�EyrVh��k^K��x`�?����:JF�:P~m8��`0��u��d�/8�a�ۨS�&@㫞���F����7��r��d�^�bҴ�!�,�3V�	!�w�
U�B!SL9��p��`��a�����i|��]���v�ߛ�P7�%�B���d�ϐ���s�A�8�c=�Y��ň�]:ģ3/�&o��0,�|�5�_�x��1h���<��+j�؅͠�,o�-��B���cC2N�B,���%�)ȅ��p�����FOv�s�:G.���I\�phYH�f2v�0��D�W�l�V��Mq�`؏ߍ$�n�/�W��>i���	�ϫ���R�?z��؜�[/�gx��ġ�v*�:ѐ�Y�k!t��B����u���l˖�h�s�5b�F�J��*ҟ�i��g|��c��ײ��Z��h~�<�<�;�����1�[�m4T83�""�h�i�'�#�{GW;�����G:�+mZ V��T�����׻]3	��ĺTZ�N�2�d"F&T�S���1��� ���r���=c��xQ��d|��i�z��hGt��Hd���V�M���l�հ���������K��C�.c�C�T��0��Yy�6R.��$����&��Bs�D�Z_��"��ڐ��)3;廉o,PS���T =�	 'L�.�k�Ǧ��:��\t�v�V�Hg/G.��ځ�&/�h��� ����J����`xQ9�F++<�xc�{��懎{�ጓ�!���=��u�ߋ�����,�Gl���CM���L�m�5G���q�m����`�Ţ6�He1A�I�6U��@p �j��/��MV���G�c����N�1�h����)%��9�no�coR]���@�xR���\��j��}޳��rW#e8����z�W=o�6�Y'�����[`N��P�x~xI�����Y]-G:O�~u�_Lm�o�Xќ�b��������	���
����P2���������\3�<#S�Jj��d�EyC{ĊwW��'K���e������(��?���V ��/]]u��v��ygy]�'���O*����q;#Qv���'���]����d�v(���g f�>��"�[�ל��!��d�l1��d[e�&�OQ�
�g[Ggm��T�(����̹~��;��cf�GO���-8��a���w��(6����_,����R�<�P�a�<��d��Qn�=�@&3�G5+}�2�B�n��Fط� @凮\\��U��!1b	8CUd��Oa�|.<<8A��o���q�(��\�:\^��>$���|]��N��qSqq��#s}�PP�x.+�b|�~3G����KA��+Z�G/w6��B�CR���&��d�}O$�Ǧ�i(�z�@��F�V�b)�'�i�C��*�������F�j"�:�!(!f@a\�1��O�) t54R�B��B��,{nB�u���3�/�t�2�gǐچ����z�@�:��=<|�k��{�SL*C��uz�l<��d��ly���y.�Oٽ�&�GL�gm��@f��p�Z�b��&a�؉K!��JʕB�\!8|MTG��-w��w�(�`rm҂�_wk���A1hb_�WP�����'��3��O�GMt����>�@����;��*f~d�g�j���P�-�Xҩ}s�M-&��@����$̠��4L�Z>����G���[������H#2f���f/܃�r)��THuH����H��<�:pzT��[���XVRd�NIm�6�Y<E5+����s�U��f���Ay';���l��H)
&����\p%��L6o��F֩����m~sd�Ќ��F��fy�ͩ�p�����͝Hڻ�޻���m��o��p��p�t� #_�?�U����������<��PU%4�>�����R��^��Q��;���[���X>�3¿R�oV��z��F/,lV6�?�Q�S��J>[_���#�N�(����nJIn��K8��	c��b���ħƉ������/$a��/M#zOҨry+�w�a�4pf��~�7��9!)��8n����S����l�8Ӷ�n6� �\:!-mA��v�T(8��4i9�dBB��QGb�b���e�.�w��kq2�}#B�b��׊�Ȓj����q�&�GB�o�e$�Y�������S[P<�Sš��9�J�����u9�n�⦾�(����<�
e�����gb-2��l'�P�5'�p|�Nڷ���]�c+���wm��
�M�1�u�;�v#�U�ț��%���.\JԦy�݇����5�%#dy�e��F����a/���>�cnǂ���>�q*��
B�,	}3���ϱ�1M9GSegɡPH�[�U�\ew:*}�Ж��� jM~��+�ά���
���P��p�Y��&�"E@>���f���1(�Y>��6Ծ���{�>���)�e�ba]��@��D�����%J�DJ�]Ҩ�����>��4�h�M 
�dL��b�.�����Z wH����;��.٫���5�|J��J�;z�c�d�l6�7g_e��0R*�3B�+(�*Q�"��Ai"s�Z�)�g��C��S��Ak�R�x��x��l�!�U"=���w�5{�����֎%��5�V�(8� ���;�=8�6l#I�f�	�s���B�|>�2. �͍�C/3i��P֒�˹�QiX������zO�cq-�++滘�~��D�)�T�`�J�������%�C� ���,�P�9�l[I�!ې���7p���)�Ȍ�&����`8���Z����n~�� [�_�
�Em��Q��<U)��Q�R��Qr"QZ��h"�Gj��.��
��0=T���h�yB�KTow���~<�QŻ���*�ʋw,�����$�;$�]^J�P�|�s�πds�X��1��>e�(����n��h0���B&�F���煄�z�'zv�k(?H;����w܆+4B��2��	�}W9��6����5�6�8�/-�9%T(%4��B��e�����N�C�^����s�	��$�r�7���R�^CL���.t�8�-�-�\S1&U��ʑ���%��3��M�`���Y]Ht�& RtS?���4�ݽ~��ZO��\c� }�eC+��\~1GŻ� ]�a\�+:9k�v��\(�`���4��֒�d�,bZ�6t�bdK��w�	I�tFW�$=���=15�0X��]/�;�eQB���V���~.:%��k�[F;�Ѥ8�5]���߸�.lt�����t�q"%�CD�CN�>�n�t��晕�`v����������e��ZFq�qpao�j@���?P�%@�S&��Âz3��d���3�ϖ�9�0Z��+\hX�(P����[�h�!��E����6�e�;n�����r��e�� 1�Op%CO�2yT���V{J8�����v�oѮ"�Rb�V�s��_�u��R�"ǋp�C�NST��Ȃ>�n�U顋,9F�%�˨[J��_�_����w� ��ø�~��!��b�����Bh�Z��|<A�@��s���b�~8,_3=Sf,���"�N�f�S����9f�-i�w��8FS.�_�xx��ۆ�.4�	f��6Au���n\%�=��;,TW��EG�L`Iɜ#)�ՂY�����.bȈ�����X����3���`s��ȩ�H�%�����ٳ5I�j_ś�]XkQ�0(+��9FaCN�T�����rm2�
ra9$[�ѺϏ�s���q�z0~N���X��&��a���SʿxBrܴo_N9 �n�	�d��J��o4,�,�17c� ��a ��� �w�D��M�;Ƣ�b��Śk鱯/s�8$_v�`���W?� �%"�/���`8�~+~
���ڤ�Ʋ�/�'"��y3�<����r8�'.�^���k��b���ˢ�~j`��"�K����F-���Y��9DB|>m�d��|#,��sG���<�?+0���)���@V�+�.��
xKV�r����ixmt,����B)���=��/]�itM>/�ɐG�$�7��7(^^}[��{�id�.wPU+�dY���]�i$��/�2r��>A�ӐA(���*��m��tòBN=����	���_�?�E���tDS��.�u=�Z@�/�ѥ�?�g!]l�-/�� ����atx�������?RQ�ߦ�<����A��;�C6�tB@���H�[��~�,D�X�4���_82���s��r-T���*T$_OI�{u^n1_$qw+y��0Ch�O��1��Y�օH�|i(��mA6�]���mif�_���N���f�RY���f���~0{.��;0��c��{c-��
��\k4����2�j�(� ��9>p�p��G4��D[6���0��K#��D�yu���?u@��J�i��V�d�n:v,�;ϫ�������@iL \���(}���Ŕ��;φ��I�s�m⠙jfw->.>����>ϫ���٢��}�>>|�	�- �P��k�4������E�� BIӝ��pZƋ=;���2=$�{��� �ẉi��M�.��Y)9��EZf#�%P�����$Q=�bc͞���\E��G3����e�^��\�c�sF� �ܲW���T@�sK~�~^�e� 4����}���n��݈o81`+� V�_�|Iu2 �ZΈ�ͭ"yI������V"��p'��	�0{��s���].�3�j⋞��y�u~��d�?��&1�		��V���+�j��m+}a��h@P��EV�7Oi��k����村S�-L�5#:��� G�E�2�FY�fl"&���W��V$zG�����u>X�gß+���dd��-q ������ͣ��p���Ķ圜 G���'��c�R�Ԇ\�"܌z�VtLk5�iV���{چTr{���Jg��B�J��o�'�ͺ*�����g���r(��`d�kvV���B
���<��,��ZYRO ��H�ʰ�����|R��}�-[G*b�{J�p"��:tw�
���Au`�L�wз恩z:Ծ�
���'�g�X6f�<�*�q���h>=�]�;��c�弳ʩ����4������`�����W�V���m L�V�sB���p�;ܦw��5�w�mWx٘e�Mߝ��4�H+�~�l�I0���?fC�ܴ�F�S]'��#��ί�gy��D��ߨ�q�g�����Ε���$N	}� �f��X���2p駫�_��Pj���ըO�cI]�����cjm�_���(n���C��'���AǱ��=x�����S�1��k�n��u�5
�k��d��i��ýNJ�,{?�����z�8ıT� �x�!�@���X*��	�lgƏ�9�n���@2X@T&�p+2b�Z��E��E��g�+8�}#�Ȩ@g�l�{̸�<A�����ʹuf
s�t���C�-S��]�W���!`�;���@\�#2	v%J-Q>��0 i7Z�j�R����\҇ќՒ�hO�>|���<��M��c�4B��Xj��	Yu��6���%��J��?���08_`QD���9j+�a��d���
ȀN[.d��OTvљ-`��o��p2X�u8	�^N�ve@�q�i�ri�%�1�H} �hցb/�6u���Rse��p��ć��v�I�E�@1�!G:	(�7zt?�i ��c�=�+/j$	�]����ʖ��gϑ)��n�796v��$b->I4����nGi�il�4N���WU�P�)]H)GW�;���'=K�HӤ9Dc˟յ��C��>����Q뙄IK��)pꑊ3m�����U#ʑ��!҆�(=V<���W,{���1u�#�+W��#ԭ#��T���@�S�s�*`���V�5�keB��{Zԕ�rK�kH�[�*��y{e{e],���p�v�)��v�ϑz�p�����a�a�Ȧ�-�T��RL�~�����C�0��P��`���<�9nd_����-��i|	@��	������{��04��~%(���W�@�m�^5���cq�� α��HF��9�sdtN��^2]q��gN �)_K����.RX�D�%C{����S��4�h+	o`���D �c.X�>lVFM����2�N+~���ч��|J�@���fE�������+����_���Q������s���^��p�������~���{%#���^篒�/u�����OL�T�9�{a��׾}XHs�L�j<[� ��-�"Ɂ$�%�GM�Ź�mp�l%�k\�г+$�.=���sF�o�q�i�����Y��[��
�����TM�����I���6�3m"���"�c&$'	�^d��D��W�R�^R�Q��$�
$�����|>k<����9��T��4Y�E�%����֠�4���.�l�Q چ�	P-���#�����\Zq��ow`8�l� X�$���|�ب@ι��^ތ�Y�\I^=� /)��C���c� �|~����p���+�dԺ��7w�<��x����8��k�␍/�Q9��i�zf�h�U��/�N��� �Ow�o�S�-����?V���:6��S���s9�`"�
��Ȧ�?��V@�\q������rG���l ��b��u�����b����!S{V��X(ן�ѾL����b!j�9�A������0��8r�{�j�Ѥ�NB�N:�$�u�%syv��
>��� �)����JF�ϖ)�!.�:>�8�f���� �}��TwA$(���?����~�]��q�h}�$���q~�T�>A�~ڐV��L����p�UR~�����w�c9�ȭ�'T �cH<t��2����q�d�@Y��2�b�n�ÆV�ъ9d�n���gCOha�AԾ~���t��2{�n¶�F��_%�*�J�o�O��.�I�gOG�	��i!lOc����x#b��A��_TF��E3�-kz�/��}���?�yTä�~_��72F5L�����z�=�J��XD���2�N�<ړ�;�F�0@ˤ��� �&g���!X�n��OT��W�6da��η�ߑ�h��a���ŭ��q�\�ӫy�U	bw�k�Nu�a�75��ٔ�DZ��x�D -}��ҭ�d,����d�Pa���?]]� ����[C>r1��1�
����~0sh�v_������BTۑ��$��|"İ�I�N<�Y�/�o�7���l_���!�#���E\��)��������f
�D��j���!����>�<q�A���uSX�ݦ��#��c��}�xCx)C��6����ዉ�����Ą��Ro� I��t�1w���[F*����������I�`T�
�G�E�t2QXr��,�(���^�L��*��,�z��N�B���k�˒���=����a�R�7u���+���H�N]�oI��Q.��N��
��Qs|��ۛ���J��l�s��g���\�@�'Mu3�h�Ê#�77IYx��&��
�0E
���ZT;��w��?�wS���XXz�:�H�UYNkm(Y+�
��.�3"a�TOd���'�~�۝�������J�u[�1����%/��1n,�v�V�;"n�z��}B��E,)-���u��rҎK2Kd7��R��A���=�x�N��T��8�Z���Ͷ��u[L���-N-*�J�XS0�Mo�C�*�$�+|櫖Y�g�S����]���Ni�r��n������%Z��wӒ��W�/�����#pWb��|�\��������w��Я������B��f'(|u�"S DN�3tz�X�`�����w��y{�o౦�N���Pw��Q�.���*��b��u��Ch}B��$��Bx����l��0c��@9��y;n.%	�OE�>��\���ˑ��S8�AZ:Tuv��p����5��1w�
�����Ƌl�(H�b_7Ҕn������&�;�u�H�V$�E���3�ڇge�rҁ.X��b�֢`k�]u*�@��N8WZ<��Җ�͔�Þ���C�1�I�I�u�OC'���ڼ;}�&�O����ԧ6����W2���/Ɲ�KMW6՚����NCv��@�I���ox:J0�|�`ȹ,fP �E��!a~_W_z���s��,r���w!�A{0�?��G�Г�o��g��Ͽn{���Ճ.LYG㸮�/��ˀ4��rř��-)�F���_�(z-��Z,8�uƮ|�eE5�XG�ɏ�M�K��-��|N�������Ssn��Λ�����e<��0@]����{��A	|�D�J�(�R��$Y���A�Q�N[�"m���󦁓�n� �l5O��VƯ仚��C�:ּ�oM�z�d���͵�Vr���jb�輩�Ob��F��&���%��,���Zi�yC&=b-
��NҝD#f��u���ڇ���k�t�c��N�}��8�Z"��ƚ�5�y�l�C�N���E��|����ޗ����T�����?s^�=;b-����0&�b���l��W�qP���q�&fuL���0egA�)�q�;���Z?���%s]A+/������rq���-U�C�4��&��#9��8����e�(��ۚ�=9n��$q.\�$�����Y�蔃O0��z�u��ތ�:/G��A�t:��������@;��I	�a������ed��YIۥ��{z�ss���ihİ�4E@O�w�AO�\U$"����K��I��M��T������[pF�g%<��>AX'��߉��X��fQ�s�}_MFґt�/-���
��\�e�~^9�����D��Q�����^Av���c�x�g�ΛU�-g?�s�4�3i��p{��r9�cg3ҧ�%�!e� ��Ibs���@�t�����#yL�İ46WR`f����Q~!�>U�@'����J��֒�[��M_��K�����5	��ᤛI�)�Ck�p�B��Q.$����ߚ�fe�&(U�o�������S�4��k���d��;�W���^~�7wt��6�l�K��qYWWX��u���Q�y���;S7x�{��������Y���<�w%熪f��&ߘ��P"���� RL���Q_U�T{F�Q��	�IE��շ'�n�#R�Q��{B4q;x��
��N���Ţ�]�Zh1y40"ֿ6&�]�D�U%.�X{��=m��*�k���Xp�#%f"��d۾�܆d}D Q�;kCGN��H',1������S|�ъb���A�A��*�C��o��\+�d���b�7)O�qJ�Y�|$���O�c�6��T��1C�{����1@x�������M��⋘�!��{5ڣ@��{_m[m��UK�bOTX9D^�@L9�ae9
��K?�O�ʟ�2$���D��	P��ORi+u��m2o�Y4�3��ߌ��ܯ��Q�̼˩m�t�;\脐����w�q��D�����?��8F�WX��{9ac�5[�	%"X#��^Z��BQ�
�7��{������4�]s���7<��+߾%	h�O�ZS[�ݠ�{�c�y�7��ew%6?�3�#�!RR��!�A�ӆ�J�&�>E1�iy~�����g������������5	�z�Z�#��n�`��������UW���Ӧ�|Of;A����{�`��4h87� ����4��"�k�k~���f�� �_���/Ә�E�y��ws��t\�O�Df�W�pmYJ*���T�ާ���83".l��<��v1*co9w��b���^{�9z��[�-��GQr�]��!�bWo��Tɽ�3S��EjhfM�2^$k�Ҽy��|Ж���\�.�ϊ�nN^����o��Κ��a���a"�C�����Ԩ�UΆ�4�5Hl�Z�O�$�-�٧�90�Ȁ*���WXU�E��&�~������_�+d�_i����~�>�toA��Va��#���h�!��{W+Tv`A�q��ih�V��M�A4�PH���O��fb�!Ϟ��).�Po�`����'����QL�"��w��Dc��ֆ�[&�:���V��ڹ�<�/J<ٿ'7�c�'��¾&����=)���`^p4s���<�JF�#l�IY���ÒY��0�N��ݵ*k�(��f&�m��"�m&>TM��\�v`�X�U�������aE�Mȧ��K4f���=Mp�C��.�1�C�����@V����V��_b��g�P> q\Х��`W����a�]��iC1A�wp>�^g�bo�A���"�gV4'TY��7�j;a�ȑ���#�9}��Tm���=A�ϼ,F86ٚ1Ȍ�,��C��=K�2C>�c��b�0Fi����j�3_�!�4C�=U\�Ch{���'{�+E^�e�MO���hh8�^ؤ��X�<r���∅&2b�R��:/C�4����<���c���B9OZ}OI	�)�����4ϋҭ��~�L֮�s?������%�	;6��sg�?X!���s(Z�f���ܢC^�������$ZE0z��3/lF͂�'ē�-�>w)��إ�����`�?���>e6*J��|~j<�9�(�`��3�y�Tż�5	���+�
�Ӝ_˜&�O���<�
<	@�p�����i\������������i���Bb�l�[�渭xk�E?ִX�=Y���ώr��������Z�Hɷ��s���>��?\}u@U�����Cꒂ���E:%�K��A@BJ�J#���tJ#)ҩt���>���?{fwg>S{f��"�]U�d���{J��ّ��ٵ���ϕ���^�a�{č(�H��u,��c�O>�i�Y�����;g���|���5��8y�@�.^r��.���5�y�9���冟Yi*c'֤���b��^,�C
D�J����k���\���:���ƭ:]μ�73oYeR8CkN��s6d�1Wfy��_�y�:d��Sq�}>;(O��eӶ���FQ6+�z�C��Do���r�l�\�~[EJШ��#]�P���<v��-���},QԒ�������?*�W}}N�7� �L��/�k���Ifa���r=�ߐ74]�+��%'���O:SF�v���"��� kƩ!
�<�����.�S�Y��z��&�'+s���/�~b�����W&�N�y���"��&1�t[\� ��{��g	'٦��Û5��ד-�@*�1��px�h5�Yޤ�ў���z+���$s*baR��|�B��<�Y&7.��E��y��WK��_�_��	+��������*���̹"U��m��)%�.y�7�.T��� [��|��@������J��+0�c�>�t�J2&rȳ�K���`mN�O��ҋ�<w��v��\_���J�
Pv����N�t8CZU��J�a����-�L������r:��#�, �˖ok��d t�����VdfSғ�*<f>���?c�"�rC��������{�[�%6��Zh��X��°�2��:�!�喯Z�(��+I�}> S�)k�.2s��L�c�1��ę	R�7���__J&o`&���o��+k�K��r��t&<|Z�����$v��GD���k��qf
:����^8}�U��m��jS���^�f�[@�� , zϙ6��Y�h������ֵ� ��H˖{������-ky)��,|���e^�|�Z_�%��ن}��o�	�XT����{�¨i�b�m�����q���\s?�ٱ�~K��*��1����q��x�Gd"FY�`����	�`��BT�]=F��7�'3����b�p!��b}G��];��m�B޻|/_�˰g�uq�!&%��wC�H���4�oVx�8���tnؐ�yx��y�5,���Y��M�z��Y���0S��T�b�������F?>A�u%���h^���nm~�v����R3���d���{�jp������� �,cQĪ��n��O1�.�E�#����~�6�}wfF����.1�;g&���y<���?����fSج����/V1�U:���.��G:X>������>�^oI���Mx{"�˾���Љ���=u�a�n}�(tALI��!|�w�s��<h�t|�;l]x���ru��<�f$�����ކ넋ll���z�J\�=�T�.����*�J��K�%U���fz��d��~�X�y��u-��g˅�kz�d}�ϭ6���w�s��T>]Rݬ�Ni_yH{������ɿOp=��G�Q�t��ryG[d\�n��>Kyu��,��)r��wl�n\p���J�fi�ތ��XՖ�-r�Đ��`L ���! AeߤБP��l��7��Lfi|�)AX��-Ҷ�g�L�8�ӣ|,�?/C3����Fp�O#P��H�ʢ��}eB���^ � L�L�� ��l��N	��5Nr���=��m"��s�Y7 >�\d�?ʶl�<ߩ�f��֩W3�	���]7�N֦u��&��@�(�Q���;�.�vV3~+���Z�i+� ��5��O��ܘf��bKXr:HI��BY��t����4z���T����˦'i�8�|�
�37aX����羬�R�7�a�}/H'��s�����О�J*�|����該��=�*��/l���I|O��ZQ|�L�ʅ�+��-�~Sv�Q�&g��H��)�}�sr?k�A<"�[��RBZk���>�N[�/	6">�X��Y�+$Z*�WJ*�T(��C�Ƽ���I������՞VgVm�/_��;����7��լ��g�����}�	���:�V��p�%䢟��K���_��'ۛn�bMJ���e]^b*��6�!��'	5\p��3|,-��dZA�S�GWp}�~���U�G�O%�2�����dd�bS�s\!bqqKq�:���m|��T����������-�,�_!�8v�\d��w�d�p��ҀO���D>w��5��
*6�c��օ7�>b#�����.����]n��[�V�m���!u_�`�.�%��#v�u����{��%�����54D!��DF�ؼ������ٝ��Q[�g���RRZs1���f�"��?=�F��VOP~�K8B�\�򎂪FR�ng�^!hSt.^&�p���~�����������Z�t��U7�*v���̾�f#�-����y�u6 �0]�n���K1q�����S���*����N��@>����HK~�������3��mpK���җa?K7��8��_����=�m�k_�A�2������X8��.�)|Wh��*r[�s@N.��V������.�hx��7=��k��G�1�D<V�y,?�f�b7���e���΄1�kv��ջ~�$�興:�P���R!��<�&��A�9Ӻ{�uZ�Vo}�"�;G	�NE��d�Xpy�5��o:�R�	x�wib*�Vp�d���na�V�(�.��j�O�L=d�qpR{��_�E�����*��˨< \��
Eq� �RBW�6��v�2r49E'n��}^/3(��CW���N8���T���#��l�0捍��	�ʬU�6�6��T���zE��fI��kA�sB06�rcB<��I��[���1�;�E���ḍcX�¶	4�8�~��RWy�4�}fJ�ź9��ơ��ݨZC>�h6�Yޟ��Z\?V�}��SǞ����\��~��" ������|��k�:���Ͼ�����w�=k�J�}^�4�NΕ��ϵ��g4�rwRJ�k݈[F۷:�<�WLR!-+X���Ǽzb��	�R}�u�/�9v�{�M	!J��ɦ�{�M�Y&Ɣ�b;A.a2�f�YTe�3сP�_Q�����h�����������=��e�ğp�B���6����L������Ul�3(fB �r�����I�jB�`i��f��C_k�d�^6��ui�=�h�ρ��Ѐ^�-�=��D0wNC!8�`R�bC�I*��� F�Iit�W0O��T���sW��+��'���m"h2ڼ�^o��l����D]�ÈMMpc�1�WDLe��7잌�8�tmF4xZ޴x��i��'��� ��Y-�!�\�^��!��D}�㙹����t�ݧ,e�5��A�=���xl� �R�{�$o��{V�q�,zt*o���7���ڔ�����ªz=�'6E>pDQ�1dS�����s�]N�׺��z!����L`��
�f����4-�)��sO��X5���X�t�VppЈ��7>��U���V��9I������sz�B���B�DS�r`+vm��"OmE����D�2#{hZ���k����TK�	������+Q����H�����x��􏮺/��j;�?�ʘ�b����U7�0W����&J������ZP'����=(������4>>-ٲ..�̘�0�M�&�%�c5F	K������c�̟�tӘ�E{Q³��	_�BS�y<锦��#��5���GgZ�|\��:��Ѻ9%� ���B���h�1���v���*�I��?�i��7y�N.�A����/؞zv<�)�<3a�f!n��syM6�͞�FK	�I�_rS�'N&�1�a0��OI�9��Ӆ����ヺjĿP��� �G�����|��]�)"�)Ȍ�E[���]�	_J�&H�\��D[?D��TA~�[F96���}��"M$��(n�dNqx�Q�i����+qK��W��h�܃��c�Vԍ[$�A��0�z3?p�\?�Zk�v5(�0%��6���U:i����&e�#� y�Ρ��D'WF��fI�!eb�����(����++�W+�ѼQ�������D���֓���p�cx�y65l w��Rk��f�L����]���?�M��K�E `5s%Ϗ��x+���E�&���~7�}Z�E���A���Fl_^�.V��8�)�^��Gɧ����W��&J�-YcL)A��=>�=b�������λ�K���oR�c�M46c�8�+!'�N���N��r����0Q�BS&���v_kF�E�;HBIFS�a�^���n���/��4���H��	qs]h�h���o�]����d@t������_�6N���C�G\���#i��H�Ӆ��,o����ʠ�E�t���G��Ե���� Q��Ս���� �N�ۍ�˦��qm���V$?��:�:gAE��6x�
?��}�7���ړHD�t��a��)�Ay�5�ݻPlp�����.�N�)0�|�2��y�%�i(��� 'ʕ��]y<F�2y:��j��Siʇkw�ǌ��a��Mw]Q>��$E-L�A�-CK��ZN&��$e��?G~~F!r�q�^�T�-~���̎�?07�`@�O,�L;H�6���:{�	�O�F�]Q2dV>��`�:����JWM�7S��*�U�N���`�{�?dG�ąl��b8t�ʭ`�)�tvZY��&�£]�S{/����U=�y�-�j}�׽���3A*�BN~9�)?w��ـ42���"9���.�8.n��ۖ^ XI3�\$���T��LΙ��*L��()v���r \�+�II��?��<�����;�-֠����pb֚��%6� ��CV#� �~�%f���X�b�{�����[������agp���D%�']�$x������K upϦ@Cv���u���h�:(���#�y�'7�|�XOZn�T����-��A�3�t��U�6۳��#Hp�o�&��(|�@��ӆ>sů��� �^�yZmJ�����k�$� Q�zt�g�:Q���=�_�pĦH��h^Bj�쪢J S�����{eb����S�i���*����i$x��Ł�Mz��k�cL����b���U���sj8����t*���%�`�>[�QOxĎohkK��3ڡ��yD���=bv1LF1���W�O9û�n"0.	�z)�c�U�u��v�-ı�����#~�BC�֛��7q�p�KRgt����-���G<-~WG��-:�oh��e�|��u�*{M"��qI��~V�3ad�iNDH�ɞd�Q�]}@�)a0��UI:q�;��9\�!5v��� �ֽ!ܕht`�388]�%�ʶ��@\|��e������(��!�����5H������X0�ڂ�%d�g��BvKt��|w���'�7YV7&Q���o�u{�I��Қ�@�!\;�B�Wkn54���ar���L^5=�t������C�l�9_CE�O��-1�ѪK��K�ڱ�T��n�]�z3�����*�~����v���PrE��e#�2�5.}R�Mm-���}_AaZ���.Y��������Y�Ve��SD��X�qQ�#���P�ј"~�?>F���^ #r�z��9�e��I0kYb'�:�7�)�dsE�w7&Į�,kp���s2��T��ŗ��'6ş��cU~.�"��I�S�b�**SB��G�Lt$H�;]���B�
Bˉ��v�>�r������R�iMB����۷ 	ׯ�2��t�F *"�I�!ܺ<�K� �"V� |
2�$��� �w�p��%�R���CMv�����J"jE�b�ď�?G1'�B�G{�0�G��#���*K��"�?���?T��6�?�M8�UH/~��59���57��Or?k��3>O6L���D���M�D�(u�(��:��fr�K:�!��V��8��R�G�]+,��i��5�3&�0Pp���<:u�1���+ }��|~y�� �j>kx�ӛ������U0���ЊɄ��&���al\�4ݰ��CƁlY�0K�����췳U��~��
���X�s�*0K�?��0�v��/M�d8��p�9�l��cjj��;��'H��ɾR#�Bh<,n�ҙ91y���s�U"���Z����GD��r��2��c�vSW���)�ΊD��:{�}c�R��F�����?�K�+�(rb�N!��a������3:[�LӾ^Ub���2訖=Qq�s�_���ya�k�N�i�/�<�?FQ�џX�N���
i�^�co����nyGA\�+#�C��K�F�7���gl�dA���cTAl�n��~5�BzB��6�"����1���ZJ�Q�V����L/�,T��ߤ_?�-�O�
�{��c�i*�\��Prv[EB�a{�ߚ!Pۭbq~�\q���w�B%�����8�A���fh��Vט��RF��Y��H��f�;�)"0f���栢������p��2�P�$�?7���C�o`@���&�B6]�<@Kc�xfI�x?�ц}}1�9U,	�$�<�u���u:>-.�L��ᣞ��|M:��1n8ls�b�<��-��R|����x����%�Jan��
�%Ww6��}�ѕ'��9���+Y�q~�:1'7���y�CH�.�`"�\�1��&`Ȩǣ*Ӻ����9���ݨ9Z�z�Q7@$�F�x����w҃��y��#��Q-�m�u~{��A�r�P�����%R��O@uafU{x|�q�5,�wqG��2l(����{/�	W^p����0l���}�Ml���e���9�5�0���X����t��]-�#z�4z�mw�L`;"w�לY[��Y� �;ZZ:%��J3[%	�����6ƕȊs�g.ފ��R;9/]t'���6�b����k�W�)�%A�}9n̃o�?P|Bi�Ơ������V�bT�-�c��WW��*����6t��3�o��IԨ��,3	嵝v�9�Y�^�^T�5�%;��Z��:��cR+p��YC2��)"R�%0�+>d�Lڥ*N&�H���
�؋�F�o��H�j+��<��7�i�͇�Ryq��,�T5������P��nIF	�_�!T�*�(U��n_,�ۥ�F�Pn(mC� �v���w�f�m�U�1��柋a�֩`�i7Ó�w^�}��=�a�i4��N/����k����!.=O`:HS����dE���m���F�0�&�Z=^w��y�����/rZ��(�7Z�M��=��Q�!ܟ��F�#�;<����gL���d�*�"�z#�g���)��E�^��|z��^�^�b��Q^̱P.�����J�ʋ���}ܻ�8��}�8��Ti�iG.����9<���Fpli����3X?���FY�aB:�����rz���!��lq��C�*e�f����e��Z�^�Xϴx11:�"$Sz�'� n��>O�*Hd��2l���<�q�<Ú+0G1RT{�-㋶z��EW-{������/Ԯ��.���blA�q{�K���S�$Ƀ�ϫu�  و�[m�io��\���Ĵ$��9��Mւ�`�$��XzM�mu���*����P�j�Y�aeBXX��b���yx�z�%%jY.���r��c�?�#�]�����-B �%�E�՗�T�<��Jxgk�
�M�L����SU�jܾ�Z� �������"�������9��4GSB7ߜA;��9�eͨ�BW˛��W92K��O��F�<���Y���cz|��?�$���Î�ý���c�]�(��i�A���}¢/a;9?藨հK��f.׸%j���3�}�F��~�� �<K�8%�B��'�7A�>��Ԥ��;��St\0wC.W��#��K�W�E��zއ�8��REq.��A�c�	���-��L<��xJ6H��]ۮU3TML�V{ź����3��f��K�0�ĔG���'���[.lR _L `���9��\�j�I��(����ӭ4)t���$q�@�a�	� ���n&��Њ~D�V��ݼ�v��e���^�e5~ݳ�~=�#t�	A�]�=	3���Cq�ى�w��7�ʻz�xD{�	��WG���nF�)F���G�L�7��\E]�p�,wG~����WL�g���ೋh"tI���N|��k���Cn��a15�P�2߰ Lτ����)�s���¼vߤ	�f7�7��+��1Y�Z˾V��𲲔���_����E��gS��P�7�l$(�Qq�|�O����� �����j`cљ�'+LO
�0�����i�8�h�sٽZ���S������|�:˧�A	��Db��hy㮅��rݗ��aj=�?�ԙ/��+IA����'6T7 i��qO�6{-�>�R�~7)�0���0��o,1��B�������\�!���#Xb��P���?Z�m���>�r��a�D?�B��x���I[1���3V�I̱�����L�&CW����8&B pW$P�r����&l�����1�)\����ѽ#!r��)�A�i�L4f���S<�MV��>ۆ}ht�V��U��	��!��zy���kS�nt�j{廰����i��a�RD[4� �'�kh�	{��Ź�/�!ʢ�<�5^��D.���@�Q��o�r��w9,�k2�\<�=�/�vIΡ�8��9��%*�������v�o�[���w�]��s��=�a_�N�G��2 ������9��.��f��S��紦��os*�>[L/�߸#��.���� ɠwݪ�A�h�g4�( ��G��
�9���I�A=�� ���\,��޲ �PV�|��D��d�_����|B�{]ks�ԟ�݄�L'�O��4�8���G�0F��zs�1��J�5"�!����҂<�_�>O+5[ǘ���{;��-�0��-"t��VDƈ��V�8,�vT��y�Df���-��z�M���K�/��k�@_����+~�|� ��[\�M��K��#F���c����j͹��1X�q_�k<�<R���%��(�&�����6�]��<+�*e�<eok�w�;��߼�Z&�H�ؤ������nW�o��KW��ܿ�j��Ĩ���@�J�i7��	簃+J�eל+�4��2��<�,�6�PYqb�1��P���	�pkB��ư��Ⱥ	k
v![���������	��NB�ѐ�ׂ�Qx�_ y�e�?H,��[s- �+l]Fc�q���/��s��(q����"��3��Q�/[t��Js��O��o~�>;�*�#}��pn�s������`�r�1܍��~	�S�������V���dO~Ò� )g�v�<��wm�[}Qv����=�E���-(��?�Ru�Xˋs~[:)u4��K"���2C�F��\��s�~��/�����	���A4��3?����8�Kwx���YN/�kl�i4Y��^p��;ia�ϥ_ �	�jҠ�G9�S�+��$e��!��۵1�h����W�C�/�&/L�͖�ʉf���q��{J0>DO�\�!+�% M����jZe���0g�`O�41��ym�T*x�kL��^��GL�s_Ȟ�������0D���^x��xk��g��#�Ñ���}cI��YN^�o2yn�E@�"K���������MM��-Od�C�A� "d�|W}�����-�W*�Q�r�� �<��.��]���Q�3�T�]au�zu��1�?s�x��0Ϳ��Lcb2X��)�gX�U�0s ~13R4�1�s��+ZĦm�e9���,�/�}��=mN<���#l*ڼI�,+�M�ٔ�h�4��g,Ѥ�5��}�y�G�i�qO���b�,���h���]r��. Sj�s3p�p/�Н�-۾{����m��7�8^������t,�oZ�e��kYP���R&6���n��9S�"��02
L�N�����kOi�e��J�U?Ȧ)��<��(
$)]�`��1D{Y,���pN�r�&lO��� �@(Ya�S'�*��1-�����|]@����=n6�riK�Ș�ڬvi+�D�m�҇�q)��&#�jvq�M�!�CN+�)bP+eN��fR���=��c�
<Ǚ����*���Grw��7��D�ќ�ww�z�P�пy!�{ӸM����*5TwH�*��iZ�#w;k�6}~'Ih�쏀�<r@NRfD�<;;!�_����?7�j�c�7����F��yۓ��/+xT�c�o�j����kZֆ�J
�k�_q��l�v=��G��͘m8`��������c�+��f7f��V=�˭E��FT�.��k��څ0�w��,����ߦ)������['�?�RV$��C��y�E�hR��h�8�$�m$�޳��a��1d�z�E�;�9j����D��H \U��m�{���v�G�����I��H";� �H�u&#7�v;�`g�ny�?��$��}��2:M�!������-�x0��HD��*/k�2�2������߻���F�h���M��
tJ0n$�W���B��w���D2�o��ҮF��?����Գ}\�\��^�8����QQ��;!��es��;��24b��XY��9�ϟ�9U';��� 8(�O���>���!��-�+:�m;a�W���\�$������oDRRgm=7:�]� ��*+a^5�Ad���IV�	�D�Jpt,��K(mԞM�^�ɂ�����}�(g��bnL3��g.��7�
������t�y�����CaV.T A�o䒼��T�a�~��:�Dl��%�Ǵ~�w�éc����C���x'�"�]�{m��f""O�
d]#�5\
�8��5�\\�+%=�y�m�fՇ[�[d����^2�X�tzr��S�w^�c�	����d,Ee>�lb���@?�|iD���>������W�O�E�b��-�yVA����}IJ��[��mz�����u=�WWNc���󵑔<�ئ�왧�Cz�A������zgU.,v�V�D���'�#�f��	E��h!5	ހ丩���C��XB����hd4�J?�����a�;'R�%iφJ���zB��-C3�M�p�����1X�9�e!H��v1���8��q����|Ko,�4����6ػ�����e�H��m �'��17�nCA\<�ҧ�����5~^3O��s]t�].��
nn�n��}U`IL�6=C?a�ᅘNLG�E��d0d`kDl�WE?��@�@�JO#꽵�ϱb`�~�M	�Pχ&�{�x��I��V
>�;GVn/�FD	LˠV^�v�q*"�߬P��R_8#٥\wiX�:;K�9=)����z���B�C��c�C���D�P~maΧ�Uy�_� ��K��Q8�j�r�����wB�,������X>�N�]�MLZ}�< �<�P����
J�>I��B�t�&[��%3����V��Nqѽ/��y2[���K���%��H��w[�'ٮ�H'W�jh����ﾼ����SUCcP�����m�W��hׅj��_�� q/�l=\�^�[�O��9!�{V�<=}���x9�Y&���p�>ۣ[�/2Fk֢^E�Э����Ah��Y@�L�O�e�t=�;��*����~\�$��C�y����Vxfc=U 5�~�� ���E;K��^������~�|ǧB��V����&�|�N����qτ�<w�̻���oj ?[o��T��X�=�G�ظ�S4��}6t����yL*j��a�OHl��|#8}��J����a#���#�lW��TK@��	*�f_�y��`����!ˋ"�h���r��Y��-��;$L�|g�>�f�t��q��Y.��ќe��5}�%�N�� -_�h�u!^��ׂ)˭��I>Y�7<�c}��|b�$!�8�(�*U��y�d�U,t��(ܣy1�q��9`�G��r�;s�����6��f���^�,a֐��k>�s'5)�n����\�]Dޟ!!ҩ����$�|���O0=��)[2��H�g	�����<t���@�Q�"*΀S!Ԥ�3�o�.�;W�F��#T�ue>AZ3%lW}�,K��t藦=���_��881ҡ�G;~D5q� ���?�職���Dy���Sk����Ib-�K45�d՟��_31i�?�;O<"�m����6a�Ju��e ���3Q��@`ɾ�}��M^��f�/�iw/2~����%��͌3��z���>vj�H�ʜcVw�g�S	�vu���V�&*q�����?J�K��CVbS3�Z�D�a�,#N�tj� �n{m9��g��������*��E��dr��y^��L���kWt���A0�/�G������m2�~��U����6*	\���&�#�7F3PB���L7G��O���q�~z0���S��>0������.5� �<|ztA?�Y��o	Ջ.��ݯ�䟤�5�\/�����ݿ��o�!�����=��_:W���վ�*�'��躿BT��j�k�'v�����kɲH���wF��y�$b��	%��ӄϕ�m.��h�������X ��Ϣ�Urg�0��w���L�g����g�P1�ޭM))�����y���m#���)�8w��ݳ��'}#fx/Sz�{�jba�BP�a5`K�2� �ˉ�\]�oa�C?:4��dYp�{�F�A��z��� *�c��}R�3l��u����"����Og���޹�{�*-K��~��^��3T�A%����Q]�7��2#���|�1\ؑ���O�u���&MK��1C̥]/Gp��Vio����zy�6Ņ���b�!�ý=Z���Q������=��N��%��"&^��X��w,)9��uF�R�T��C>��,|ks|�$e��Fw�CC$!i����ы��1;���f�ŧ_�����^����`'�����X.;��mh���TU���f�S��)���+�ǚqٓI���6|�Mk�)tGбx^��CP�#�nTҽu���'��&��4v�v�N�v��Ad�!��ax�ad�ad������D�m���*�A�/�נz)J�'�'��sf"��$�m���a@@<Jd�I���݋���^�P�}�ܳ�?�����/:m�;w	�m	;?��!���=Z�2JT�k�L_��K��;j��St�Y������mtL�fz�h��8I��N����OM����2�M�)��"���'���vH9�d�y+�7	��c_�G6q���.���3���fa$�7�Q�M�-���SZ��Ew�����jO�x�$Nb=(���?��,����ZΩ�'˂O"<�Y5�*cC(��mf�:�f�z9�Eve��L�W%����_�M&�6�U�fX�E��ms���k�[^�z(���u3��.��~��.�ɨ�!��������r�M+,V��7����O�#���o�CQo�z&4D��?y�t���b7\	���c��;�ja]c�T% !9
�eG*���`#o���W�{/��f�4�lm�*��-��������2D���*��]��y �g�a��R�b��Oc�|�_&�^K������ �KF$�iF}�јA�����Un#��u�"�&��ήV��'�O#a��'I��k��
�ۼR�c(E}�9�[n�~��m��ӺL5�,��+� P,�M���`����H�R�07>�8��x��Ѹ�� ��,̗B��oo�M|���j eiK𡹃���	�_u���[�u�>م}���I�[6��n��|��A�R��*2~�����?l����s��O��!��>�o�+uh�"�(�@S�Q�ͅ��ᓺ�K�1�#���������QB�$�J�����W��o�7�����no6���{����}���{�5h����d��4k�x�u����Hh��Px�id,(�i��?�i;)��9��A\v)����,7\*���S���<����)�9�����zv����[�5¸�ƮgɕG1�([��)W�^�"D1�%<�&����_��|B�Tu-���zBx���������T,8���V���C���,�8|w�TdL�D�5"�$��Z�*�B�z�&���.�w�Y��9#O(Aq�'�qf�e]�;���W�]:�	��?��#��_b��1Sʨ�Js�"�N��b����
aW����t��tw���r�'2��3_���=�ye�M�&����Q,C
=kyR�]|�u���ݢ�j�����<B�ǡ����lVua������5Y;<�EPC��πn��A��?��.nk��P_�a*�!��R?����
���0\cŷ��Y�5/lj�j�;�P�@���/���Z��&d����pꮟ����?}~KT��C�_}�w��lƝ�gV�J�h�{��r��نP1��p�Gq���/�V#%`$�`��겔���ߴ��*�ɻF�d�󳍍���u�2082��?\�"-S/�j�չ�+�t�ޥo�4\������j�w���
O�������
d,"�D*���3�2Ǟh���P�c��H��hڦ�ӈ�����!���v/�v�B߳r�(_��!�'���N��!����҂����i]V���ݛ��؈��Ki��>!�� ����J`��F��n�7�@��R]N�6]��a`1���BV"�T���U7���(QϽ\�e+� ��ِ�ֲ#��~�C�?���?�[�=���a��%")��1(qz�.��x	1zny�?o��}V+��K\M>k�h+V�I����pwW御�4���Ӣ�;1�
R�F�.X�vj����8�Y����㓄�b����������F�0��<�'��_+�Nw��K�oh�i�]~���;;��P;Y�n(^�9V�h��(�g���n^��~\��T}����7��wд�k�m�(��E\g��y��ܴvU�WI����/�<�<W����/�	��ӣ�����T�Ry8g0�G�'4ӟ���PQ�"~�+�OUz��hsC��� AU�/u�ڸu����F�*��������gO���o��C֜8|�*���T#~,(*�2u麇���8I�	0ή�*܈~]���dxg�(�TV��Gl���� ���u��fJ����@h������M���*Ù\<��A'�T����$/]Y�`�]*4��['�j�2:�>�z��ujp_����tf�gJ�p�3�������o�$��r4�ɨ a)���R���k�U���4�wު>��"n��-�~	V��S�5�{9�m�S��~n�����(����ȠqaIl�i!x�A|��>��Rpk'�� ��b��y�KI�Ͱ;�^�ji�g�9��}C�1?�IS����+�60@�ʖ:�(����rx1zӾ!�^(�w��ΧԸ��b��S@�pr����)�t�� K������3�Ԭz;o�OI'�{�3���妍�
�ӓ8CK��3�u>cʔ�s7:W��.ۯ4g)���%b�N6k��K��{N�������d~E��{��Ln:=%d��8[1=
K�ME����;	�_�Ǹh�ե��OP���'��A���ꦲ���4И��ث�O�>�a��0y_�d���0�e��9���!��}!�ST�/f�RU ��X�'�ͧ{J��/AG*�~�ŕ��!̲ٴ�L��V.,�N����`���� ���P���X��x�N�A�M�J���'��i_��}%��C���D��{Q���d��K��/Z���%؟�M��yex��5���.a��߲�~��$��6
������.��KS�G^��W�?�K�>�~���=��ۑ��a,�r����~2{���	_X�0�P��NA����	�1��8�O�g�4�_p�zJ��Ǔ�������Ԭ\��i?�bZ��S���K\E��U�n�L�擈�����x��=�H�M��\m�~���@~`��Õ�g�i�_�"�V�L�����r��m�����=)v�����H�q;Ӭ	�~
>�=A��57Τ����:�'o�1HU�-< Z%��z���%۾�Й�- BX�QY�їP/�K%�gj���O �I�`���g9�` R�x��A��"�L��{�	M��0��Tx����s΄=.Q�T+�f��P������F��w��ĶRZ��n>
Ǜ�G$<%�
��U?J����bT����(�isM��o��~��}���*��4L&� ��)f��#$/�]�H�s�}1���ӓ��y�9�x��6y�_5{D��'c�!�;�mb����nɖ����`��M���rM�]L�����<(Ȁ��1���������~����K�b��M��V��)���L�ȔDI�xG,+��8��>�N��4:���^I�Zo�G���T�Q\[p�5Ӟ|��>�����<)H�1h�?��t�P���^�V�)>>38�/�<���WV�z��"�V���ͫ�E�*y�xʀ3`?\��r�	?�#���ؘ�|�&�ql�0_��ȳ�)�͐3�=��\=�����f������'�5r�8�p*e��&���WM&3���n4�ƥ��=��EU]���:���i�3�Iy� �Z��7F�gH�	؏+��2�̾cbl�e?�%�hu�6���rA���6�5��."ؠ�/n�\���ٳ����y���ޏ~�e��m�f8^�����%W�uTI�
�2��|��d�W�7���Q#�B����W�vӉ����9��--�)�։ w�٦ݥ|�����&��S��*
�<r��4���,ɣ�+`J�7�	L�"��>�^�����r>ǵ.[�X���Ѝ�D��XJ��k4�Mo���˓��C�G��� ���վs���>맜��Ǎ��x�ݞ�gyx�G�<�;�k�>$fؗ���-�	>��G�������c��Qн��x�hx�n���z�[���祵?}4st"Gi^ƿ����>�Ęn�!<*�i���ѱ4�D����G]�EIJ�7�-���k�`��^�U�K#�t�
J�4J� (�݈ HHI(")��]C�
�%�3�0���=#���_n}����ٱ�Z�X�\/lY(��7�O�|�FZA.;�w��$��e�QwV�"�� ڑ����F'hL��u�TWU�{�s�+��qG-����t�g/AަJ�	�T|O��g:���Ay�,)�(�����ܿ���
HF୽��_E��p���R�j���O_R�OT���g��>���1g���ݜ�9�\�I�� �e�������-P5�!����s���R1�c{&�r2:M*�������2��h�����C~�?��&Z7��E�m��)��>>	OoU7���Fg��*U�/|���yn?	r���G ���c���/�Xј��zU�Ϭ�2��a]Ef��F^@��W��is�W��Miz�s+��lB�.����cSF�z%=n���CR�An�����[��nug����]X��F��dy�F3|����1�.B���1j�������nW�%Ⱦ�iZ�9�y��>�^_A���[������דe��V]H��X�t|��ZE��Kq�dp������iⅦ�,�)�!S�U��@�5��8�F�CT�m�r��,���,��?�b�gb�ˎ�.)D݃�l�_O�Y	��%WO�1�\��BD������f֊�Ņ�/�e���Ҵf +��O�4����k~�:D����Cʫ����W)�\*EU��\��D�j�&|�]���KMy�͔��m�{�1*��˗�e$��;]�qmU�alg3Uݱ��,~A��5�vp�����Q�e+_#�pc,�/Z5������5J}[M�<��y��x�OF��\6U(�:����E.�')VV{�K������M�S ��iva���!�o"G��@��YF��O\o��������nq!���P̐ʕ.��\4+ox-��(B�~;��˄�}` \U[����k�TEI��y��ˀ|������77�#pdJ'�Dͤx���K��ROFCYdFy��!c�I����\�PI�:A,bqٌ�ht]eM�'ϭq]I��٩\�q�Gj;\�՞��Jѻ�=?�"��+�����v�"���~yC���U G��=dK��.2�����1B��~D��{�U���'����,#!3�Ճ*�����rt�\Ԇ`ݻ� Zm#�@R�
�0[�_�?��J�.��Qj��e����A�:9(��db��]�u�<�-}iyp����&6�?b��YM�: +��G���wD/b�r�Ju�s~sͷ
�'�2oq���L�5��e��L}��F���8d������q?����.�#�����6�������Mu۹���_�>�f;��h} '5�y�*��*����������H��_������n��
����lw�w��7��	3��6��i}��k�2O�3e�u���N�����:����"m�vI ��Nu�7����w�s�L���)��C�V�PB��[^yr)˗X��zO�&Ȍ,��U,����p�z=��չ��NÞp�rd�i`-S9����^Ď���r�aVS�!s5��4�����,~����i��wK�eR`� ]���\��ت�^y�L�E�õ������ �z=-�z\��aP��iH�� �\�U�1���ׂ������S��S&��531��ĕ9���ޟ������z"�2���Mv���U��G���Ow�~U�Bۑ���4K��D�/|�hj�]������g���a�����/���a�}{�O[OI��g-��s{T���g�nʴ�y�Z��^�&:��ͱ�Q���+c���[z=!mw�𛿱1�-����T���&+�,"F�t�3���Z2odo4�j��F��ӄ�XxD�����p��͂�i�Wp��W��� �F6^)����c��w���	��$@��}�1(3��7Yf@m��trr��ڲO�+�/��ZrOW��H�r��?][��j��+;�q�y����g�E/saG����/��_L}�Q�Cit��c���S��T�����`!�4ѽ��}�l-���u�Y�pB���]8=��>|��a��ͥ����}��gH��1A�W��A,vֆGG ��<˞��l��6���т.�+��yջ���w�[� h�/�U����⫧sn�N�M�ʛ6R�ͻ93���߮H��z��_̿�2Jس]��`��s<d�sW��3������9Y��ֹ�M9�����L�ҋ�x��� �C���γ��]�����I���9��R���j�@ʗ�Fgǃ�J
33}��s�z
�����k��8�z?g777L�455O�p�3���"��I��)E���k��F���F�L !�`��@/�L��WUUV8�z���8�C�����#� ������$�Ȅ�@Y8�7�k�$��dS��p��[ �}���L��:�U@���%�� \�OL���Y-E�����\�ę�,��:�� H����7jr}�@�]��ۇ��>��!���&��f?]3.@+m�n-3�,���-�4\�[���B���&U�Lc`��"A��h'��JS�SE=�y��'A�:�T�?������~������s�X���>����Ʈg[�E48�Z��`���ÍWq��H��W�����`���x��V˕J�}�N�9�Mo�	��%Gx��)�ռ��(��3+`O��Ҫ���]M�Ϣ~��Z}�y�<&p5������/fT�0��ߣ�|��99�z\N����X�X�u�I�gx��2���_����z���]��8��<<c�*_��5���թ�`,�� ��~B��Y i+��[�b����@������}!�S�0=��h��D�)�0���׎��A�3|��SԵE~�<��_K<^�D^��`�����C��
���$;�fϚµ����}ĽN���K�.��g�$���6��V���q���s���t0�W��Q��g^�4�&��a���r���3��i��ڴ|�1��x"�64^X���m��ϐ&>`�j�=��x����jLC�WCz��Q�D�v1�-���ũ�kG���wvvN�:� � CZ ���fE�X��|#�3��X<�k[=�����k�ͧ_�D\�����?O��x8/�JN��0�N~�;�ڝ��[��ɣ��Eq��)-������8f��<@p�| H\QQ�@J`����@�l@�>	-o�� 1�i�H{��4�X�;��UYt��x퇀Q�K�9(6��������q�����;H�L��*�Xz��LMna!WsK��yFX�<6?L���E�����2I��T�!�@�y`d
T��:ո��kl��p)dɥ��M{/��f��[Vѓ��Ǆ�����jhX틭��~���y�~�+�T_,5/>V
3p�Ó�����rw3�z���m~Y"k��֝gg?��{A�k���wW'QF��!���W�+ͻ��Nm���ߺ'Ҍ~��)#Ԅ�52��~0��R����Ih{��X������x:�ڲt媤$�:�����PB�x+��KN��
Rͫl�.V2�GL���|´�9w�YA�m��@ʭ�D�����a�?\�[�2���?o$�5��l�>�)0n3��h?���:��.��o�(m��hw�)��P�G	@��~��^f/K&��8oc�b��=��V6F^� A��^���1 
@�[�/�uD��|���G&���g��K==����� oaa`�oS���8�Rt��?HO����3s�Jmߤ�`a&`ΐ159���mx����lfB�fMol���f�L�3��:�����:##��j��L3�O�3��TJ��G q��1eg�6��(�����t�K)���{8&Wmm�_/@�;D
��J{9��dq���ބ�[������v����?a�8n�qo+u�M��T�Bn�y ��o������un.Մ�5..�S-�jF=$止[|ǔKݻ�7:�i�5�@����Mc������������7H�O+�*��Y��ζn��:;O4�&�$�P弘PŢ�H^e5y.��(����g��s�,O�&m�pn�5�,.���s�3n���J�%[��R�2���kz~�شl�8��Ē��h֦�v��Cֺ���~�Z���KRc���N��Q�0�u�������v�U��^H�e-n�	�oxJ���^sm��rrTd����M�g���6Y�W��!��5c�����H:
8�q�b̈�3�1�<i�_�mEf[�-n�O����ɹ��f��� غ���y�
�A�*�����Z���H8�R�҆4`�3�v+!�8�M�|9���,�"P�W�Ld�ᒕk�\�10hZ21�r�X�)��/rq
|����h˰ޯ�´B�m/�����"�)���.�KY�;���G,#�N��V}wd�
����~ʂȝW�_�FX��G9ۿ{�I�RGD�Q�A���X_�r�$�̥ԫlJY����|�r|p�Q?�hU��u��C�i\򳑫��*�L�!?h�U\�O���m,,sm��q���J��E����ҾK��Its�#����lW/��1�8�������?P�y���M�2]-��s�nӬ7���>�̽W�gNa�/O9���m]ʠ����������%ޤ��z�;� �ޅ��Y��v�+�G�I[
<�b19(ʴ�nwC�m�R�c�'C�;D#���3J��B�cY|��o�ʋS��f��ϛ������3y-�OieE>��L$�юz~�{aO�*h^���-�r8�+K��0g\g�|A ��/�� ��K7�� � �>���mh�b���� ����x.��E#�k�>CR��t0ا��Sʮ�`F'q�-��?El��R[�>��]�*��΍~�d�[�	C��x"B>���,�����6��H
GI�5���O��}*~���<�q���#�[�,9q�r�K�nd|������@�����K]?l%���R�Z�*'�*�^f=�����5���)Y^����?�\k��߷��T9��q���P�:O߂��d���"9s��?)Z�~B�Uvϟ�N�6��	�&��2�w���v�r�/��*�9�X#�&r=Th.l��8D�,]�d���y6X�֢�Gu��T�ȁ�H� ��ʯ�p�"���)�Y�^�j�^�.j���st��o�	De���S�������4�mVr�.�B4������N.�=�Uu�ߛ�����k�`�6��? ��uD�P�j���B�em��.�T�3b�ghIRjv��n00�
��wH#��i��s �Q�j?k��%�V�(�����#Qtm��ǝE�W-�4��JETĎ�ϼ���Vg�Y1ί_G@����Yml#^9e�3oT�c�
2�Ł,�����J;9�3�hE�] 9wO�~���f�*s�b������<�W�����ͦ���~��

�d5V�E�iv�hme%�	fP�"pe�|��gqŶu�E���>��Q]E�$����Gn��BaV��� ��R�6���ry"b�%�yl �P�t�-/sD�:;۽"7�ZX����Yj�k1�����4*�T"M��P�wZ� K�b�\�j]��!aΈ�ð�Ŕ�*��a?������~<<_rdPN���K+d��"X���Om��-��?9���ӹǛ%(We��9;Q/����DR^�Ŗo�*�i}5�U����|��H��o~�P>��5r��j���X�`�gzX�X����{?�����#���w�J���h������z�c��}�n�{\s�B�t&�Cs:����j�3�'i���)dA�o|�0����GDaM�'�>R���l�M��̉�[^�j��8#M:9�T�����P�Dٝ�>����#����{�!0?�bv:z���(��3p���X�kR��E��ww0w���G0ݠ���z?c�|냜q1�h 4�66T���#Ng�A��l	�u�ϒ���>��`䂆/'�%����t�k�����3�=�ޅd�=��4׸>���6kP��
��}�y�n�g�g���0w�0�{�}�I
�����XX[J��J|i�c�=�SI�O�ђD����^��k$`o%i���'�<�(*-_W��K��� y��aE�������9�?'[��NF�$�A�J��*eB� K��x%�>�y���msP|:yǁ��૥��f)1��>�~�c�i�^�ت&���	ϫg�Az)�v-�@��T�Ydz���<C� IFW�[��䠵R�%���\����i��߭I�/7a��PH|����]���g;J��T6�t�O�n'��"��/E����>�Xճ%'r�i|7�|��_Y4���PT�%nc��
���S>,�C챩bM�L������@Õ}�eM�/�i>��%�$ �3}�#��o�m$5�����<9��9ڱΞ���S��M��^��]����*,%i��vs ���~g,  9�����f�b�b	{�٫�"�E,b����[�R� :U�ٺ�疯o�9�H�����N�S!�T�w�����W���>&����w|��Sd��Ծ8��Mc��l-
��
� �%2�WY�ygb�T#*�0��l�{8�G`��H̑���3$����
`��2�<���z*�+� 䂓 P��ް/?��btJ2�	������.�"�ڀ�bҬ(��4�m��F��d3�Cy?�j�NF�f��O��Q-ЛZ�}B�#��L���޼
�5�i#n}�҆�:�CښPh���ȣ�L�|\��:��(�Jv�[Z���g��v��)c:xiy�,>��<6�W�P�$Gp�B�(Uu���/�ǧ�XOe׸�af�O��6������k.
��}
Ծa�\=�pL*�����=1W:������$D�ʣ/lxr��nk�����'�yhs/O
]�[��ޭȤ�E�Pw��i�}�/�1��_�0��0�U>{��@V�8�l:�s��M��?<���H��B'w��&3��HĢ�w:�m2�t��u����L�Ibn��3[�gKy�����:9H�%@� �Mo�/9�s�L-Q��ܙ�T�J�=J���8�}�}��T�����'_H�Iu�RB�����}>4� ���D+pG'�2�	��yR� hQ�������x�g�I��#؈j�` o�����y�4�,w��������Uin��� �1{����"��/��%�@f��|�_�N�҃�;��g��|�G>�8>���C,�����7����\�S�	��Qi^v�[�ۯ|��lu��,��n'N��T����f��f���_�SaIĢG��ʖܑ�I��#�������SG��^�]r?��|��}�{�
]�����s�z��%(��/Z�ο�mݴl�JӮ��y,BZM�|�����k�����O~Y�}�ĥ|���E���ј"->�Ҧ�m��)l���,���?7#b����]��'�h}�~���{AqmNB�x�_bҤ*O��?�Lp����NV�}_�{�(����r��dȜ��џU$�gvg�nڏq�Ѿ�퓲���xji��u���	qYA ��3���X�����;��^Q��>� 	:h��Y�Q���Q3��b���Ё��NI�rIx;�EX��g���+�0v��~���}���,�5CL�;���?[ �Ҧ�m9�>��8�A핞�7N�oR����z� FXK\f4[���l��u5��3�T2n�c1�!������įDwE��Y6�"!h��-<q����#9��{�j��Z���$t����!��օճv_*}Y����'M��X�L��WS�����
kB�A1�7H����9:6�bW�<�o"h��CN6_�y�=ZH�k"��vG��R��v8�]W\;z�Z�U��ǩ��7��&Χ�'J�$��\�\z2Z����6�+���L��G���6��f��C�DY��R�?{��,r
�`K��a,�V��b"�S	?��+�-�+k�� [3ȸ���������,[���u�7rЗ�8|V�����{���r�o����W��Y͜���X2�����%�uG&i)ԙ���B���R	>�|��4e�T]�B4w�q 9��lX
KL��G���
_���e�r�8'tU�Hye�o�ZDWz��h��v ֑x����	��>�i�X�@#��&�J�+K���r���a�<#����J Z��Z��JX�k�*�}�&������dnr`��;K�52���ƺ):���˛|��.LuJ��u�Uz#�M��=�cڹR���L�Tx-�O�~���|#; KA�"?��
��^L���3��L�f`�]dy�L{�M
6��v$��H`��BE�f������H.T��L��ݚ��c�奨Xp����.1ќ-�l#�	DX[�_�w%�K��"��|s20�~I�(m��v���������h�����^!#2�*Y�V� #�3���H������c<~���	��Ġep�)/DKRr����Y
k �=+J�J�t���[�h.wH{������	ͮ�e!����-�U�L��Ż�ݞ kP�eޚ��fYe��.�"���O��XFv�����L7�A�lC\����H�����-��O��+Me�� ����rN�g�¤��N�;��$o�˚`�R�Tʎ\��:�����iO�}�w��+Ow\�T^�D8r��֬�9�_�u��Ӵ��p� ����ך�]�Ybs�H��s��U����~���lg,q�ʣeZ�%}��W�1a[+Z�A���Z����)���f��iQ�R˻��v��'*���r,ؤo�5�Z������k;"M��X��e�U0K1�>��|HNĬ�3�^G�3��[�5��1��ŉOP��e�}���7��5~X�lI�3�Y����X��$ʡ��]s��la��`���W�d�0���&"w�Mv�wI��p;a��+��1�����97�s�iu'!�Y ����.ñS��������fQ��	+H(�O:�?�Ӱ���B{���]. 9?�y�!L�l��jK�pɗ%�P@���������6���KU6�s�?���,��9+]qi�]v7��Z6H�|��ǔZEz�S��jI������t�cRrԚ���|Ź�X��܀�h������*d+��Z��ʾ�(F`T���69�j��t\�A�!�E��T�[���'-T��\D�t���-/�&@9�̴`�^��V+���R�� �����Q���ƖP�?��b0��əb��;E����#
��Q9�G�e���O�K!-W�)�6L��%����������|+w�N����Jg�A�R	k}�}�hۃ!1
��b�,����O�sdE-O	Z9��h`�����Y��3b N:t�{����"&��j�78�[9~�_�o]� iG}��#�(�k�Y.^�%6��)��o�����fM��_����'����6����
�7�� ی)���"��K@�CSS3+�`ϕ;y�����k8��~կ�-��ꝊŅX��u&�˃�e�6�~�*`|�B�΋'���,�g���z"�v�X�$�O,�m���
s���pڏM�W7��ar�Aؠ������U�"����p5�bz�.�����"��r%XݮEK��-s��Ӯ�g���C?&�D��V�|!c����b�UP����I���f|h�孵1�����y񋸫�;��fM8��O�5�7Q&<�O��$%�;�z=Q�ez�p
���Q:.� ��:U;+	�Km=)D��9^�Q$����۹�Kr�8�	k�S��t��5�md�&�z��A��;�5�(TҳP$	�`#�6�J�n$�y�R�4|
�j���e$�8p����TQ�淌�?��D4��fw�޽TKV��|&�O�&9n߂eXO����$Uw��Pi_�T(�Ҿx�葖N8�[�}r�,����q����x�y��hA6���dЍ�_ћ�%WXe�'�����5��c��P��f�A�#RAR�L
�&
��#�(8x��Kم�J� 
��tk���(Op/W�11�j�g1���9�y�����Ac`�G���k8Z������ɂ�g
/��F�Y�������X0B6E�*ƣ��l�#�A��N�oY;W�cNn<Q��_m<%s�f7*z�T�3*��b8�SQ�o�A����.+SZJ���$�{�]i"�ͺ� �Xw�C�gF4Y��L�R�B�?��Pз��ի�Q�����"9x�.���;�����Eę�R�;���xM�v���@^�Z%Eg���\@"�scij����A�����]n�\�R˃�HE�,֙�;��Wޞ�sA�t�<�{��t�vh�[`]cu�����0$��w2p���_r"���~�3��@�A�8(��T N��-�7�v�>o��=�ZD�9@����H��?�r�J�p��c��b��Ə����������m�V�@�%:saz/�?��v��,�e����=O��ҾY�E�8�2������:��ވ�1����e;�<�&�]��k�g�j6k��o�Ȼ=Z��[�����ԫ(A1&�6Yv��_~���q��(q	����zl�/m�.b�'C��Ǯs�h��R���h.����+2��ߏ�<N�姈u6;����(Yc����)�dY������X�$��??��� �c%����Y$K�·Q�����0�y�}�y֞����l����+.8�G��حd3̎�aa{Xق�Qk����H��v���&��!�lK�h�7?ή������������ſC�G�܁�2I��H��h�pC 7��+��u�a�6xX��x2�m'Z���WC�O�H�V6�����z��@�)���������<�i ��9t�"c�zO|��-oVE΃v&^�|{�c������f7؜
����?8�տ|�o�
ؽ+c+61��l���{Q��$�l��Z�g�,B Y+=�X�N�a�>�x�TZ#w�2*�@����b�S�o'"V�{>S�������Q�ءZ!�9@w����x�*'�}�aMV}Y���8]6!���ŗ/��X����`�������]%��K�1�T�E 2r+���]Β�a�Є�x�]?�8*Dȥ�cw��
�J���X*�k�� �OE�wr`[�a���FE�Wx�g���5��FX(&Mw�r�&���t�
�?B�4��o8/���e�@�d�|��'���Rf� ����
JT��X�L.#6[���=���=�_�ìv�R���}IX�� 
)G`:0��/+a����\鷈�R���y��D�@Q�81�n�_N�cp�g{,d�Zᩐ�>Q�+	���C�;f��~�-#ώ?xN���} _�˱R�~`��:�7��bFg�v�B��
f��'Cᑦk1�k>�!�v|x�l(�T'���Q�L����N�����*��d�xq��ɿ+����U�1F�\��m~�P�=�ڗ�?��w+ "�ޓ�����R��"�j*K�[@���#�^afgXΛ�Lb��h^ܰf��� r����R�&"_��a����)��JGk�&��d��g��u�I����@�r|nRa�@e Wu",�k�������$O^�ڮ���Û�u�Y&&Y��I@���b;���c�R�h��y��>�~�P��2��v[�Td����ѷ2#�M�*
���P�����UϗY�kʛ�k��8��u�{m�~$g�r��T`g�ѭI.�@��_��'�Iz̼#$�@:�5J���/)i�Q�e�.�司{�s��<:��XN�� -�߬����$o���M����mN����~S���'�&H�{$����pG���x.a�DI�F SbN��{uy�C#�Ng��dJ����3ɂ^�.JݰEv,,�b�<}NTjֿ[a_`�%,���&�3�:�����*�Y���@�_�i�ݺ�&sN#�1"����kq����H�&�mA��Z;�vU?���}�>(K�ڻ,M6i�����iKߐw��e�,`��i�|���1�F051} 7�g z�?O{E�����M��]������r���͘ҹ�~�9�H(l��2q��8��|��������@�t�g"S�dm���Gз�r�w�z�X��*�q�v�/�#��%Ȼ���L�Q�v�>֧������ t��c,.�gA�}Ȏx�ލ�uJ�{�W��U��a��/��W���$td:?��#��:e��1f�r��ؑ#�u[�GK����v�*�d�Ĕ)I�B�>W|p�/2:.W�{�u��2��8�H���v���:��-H��B��������I����x�(!�
:LA��z�>��<�e���&�s��������� �l�a�'nM�ܬj�W�5�	�	@B�Bz~��;��C#�8�J��YD[�*�W$���������0\�ή�m�#
Qd'���P��t�[K��_)�N�%�1��O�PZ��� HsEQ�#��'|ҳ�t�����u�@����t�[[�F�M��;�(�:y����Ԃh�S��KS��������Lj��[s�+/ ��"����5"� �n��\4�?_���hԑ��2�+�WMW��wW��;�yk�aRz�y�%W�t}�F�n4?�PT'�a��k�*�E����j�'�O�I�!1��@�xeQ~�Y���&FR�P�ϓ�cC���]�')������������!�5���c�5\���y(�k{��;$�NCl��u����#�Жp��dA��0>m���#�ۿ�D(����R�	l�bIZ�Y�?��h��l�מ��N�F�S�w�!P��sgλ���I�������
z��P����������B���[��$�*��RfOo�$vO4s�d�{��[�L���}R>�X�����{!��k�{�#��4�Y���Y���/���eVs�"��⣧�P�u�bs[��͇��j��Gn���#��DC��y���!�y�aH����hJ�L�r�h�1u��,r8K�UD���!�)�w��X����l��B>��1�u+A��D����N�$���Φ�3���bSt�x�p)�z:G�;7_�䋫�i�}�J��=�WV��ڣa��5!�Q�7R�Y���JX���S���Vux��-B�n�L)�.?'lՐ����XQo��ЩRߙ��p�/`���3܂)lPp��	4����q�S��L�
�/�T���O�.��P��Gʂ���
(�]�ϹO_*f����F)���Johԯ����xb��n!w`A�N�R�XlX��F|��5u��:X@��E*���0E�U�$�T[��>o�ԝC�	���_�� fN��r:=�ƎrWГ�(*:�V�~�ϱ�Z�T5�T�
��~q&I���ؿ�a�M�ޚ	 �(�������?�+k�B��<���jG9z���]�'4�:�e�$�ⶱ+FwT������$�-d*#��D�X�R)!��C��rC��I/h ��;*�f�ۨἙ@��Zfr-˶zFH�H������S�P�4�}�xc��[@��:fg�zU�-�爏��P�&}崼3N]���y&ҭӷ�i�?F],_0��Q]�o�؍�/5x!b�u���S�ς���׎fOE$.�?��~�]�ӑ�߯[/�S>-I |l�����_j���pͲ� ��4���#�T��3.�9�9_��@�/�i��{x2:�5���p���c z���Ѕ�l{^7,4���z�v��J�in*y�A�ǈl��d����֕�}i���㍆ϐU�
*{��z��`iK9
�m�o�Z�ą�fs�W����E��������x����S
�yһSV[)S:�M� =$����<���L���Z�r���dg��b(�U����ڞ��٭ܝ_yo+��b|(�ܛ�QUfu�������JN�`�gqFm���Jzv�7��n}���K-4X�Z��6c>0+64���Ҍ~Y!��s�tb�	�L���#�y7�(wD�y�8���sYLy��+�J+r�.2io�
��-\n�h�i����T����M���*��+Q�Að�WP�V��&�si؋6�3�AbrTRbFlGE˫�-�s*<�z�)g;L��Mv\؛�ARP"�	�{�,?��v�>�ɶ
g����y�;$G9�r�����D�'\��ә�Uz��L!����r?Z��;,Cs�.�q�Q���ۊs���
?~���A�}]�F�y\)����L�٭�����B@?�^����w�t$L�Iu#�����������0�������
Je���8�8��$�N`���D��Ū�å��K.�w/�T{��K/�S��&^�\_��圿:M�8��ԩ
.�j5c<���7��,���ދs�ro��7��3<���]�' ������dCb�&}�R�۩`�?�HKP��x�A*"��HS��Ty_��o��8xw1/�p9��M&}\Lj����{
�m�Q�l��,��A�C�\��ᗈ/�Q��	��<������T���e�Y���6N�d`<��u˼�i�~�����b�l��2l8�����PTb���քxk0���LSsarS���Y|Bk�W�a>��F�|w��� 1���qS������߭ZG��G�F-U0�V��Ń�l���ùX��K�Ҵ��Eq%V:���jߧ����+>�@���{���IϤ;N�_��G?��x��ԟm�NJf��I<�� 5˯�e�~���������>�;�?��I�q�����H�"J_�Ł��vގ��ſ~�r���X"����w�0������ºe^�A9Uݲ�a�w9�Q�K�br~jD�~�Q����v\��d�˪���t�F}��+�c��\�|)�Ŷ���f����|�����Q8�TO"���I|�p�<��G����H�E
:&���&��?�^U8�O�z^�9>�>M��Nv�u�e�=K��(SH���5d�p:6_�v i�O^���X,A�baIj�b�g�?���ө�<'t��L�H/K��(��' :E����7v%�+��ܘunPYr�~6kq�ᢿIݷb��{vj�>�6���Xllw�A��� �m쎠��GM_'��?�_?���{]g_������+	�u���0����	$�zSiA�	��X�`�sYX+�ǯs�Ϥ~ w��a^��<�I�%�p��7��Yi#MS��$k��ޗ��5���?�����n;a2�111qc���#9s(���;;��%f]jW ���ܥ����e�|����>�f��]�S�Į���N8>*�����y��4��>2�I3�Q~O)P+.�P����%
�E?����ӵ�"� ߗ�,��g~N�uq,D�?'�m�Tnl3Y5G'��o].�j����w�b.G�fҖ�����çm@���P������ӡ��{N@��[eMM�Bڎ^�,��3����]���·e*|�s^#e^�m(e����"���"]T_wz�4[�L�܁���߈+D�<#���x�H9�4��:���$|����ݳ�Ҹ�<��o3O��K�E�ۍ1[f��g��Z�&oTnϸ<�T��cU���N�W�x���J���8V
'בQb<nV7c��lfKLm��{Ă��F��V���'�͞��W�O�oI�Rԓn�$��5���ӞFY�>��	��y2��d5c����b=��s�]E��e���������byY屮a�4���6P��%ft =�){b *�_��:{�⭣]����U�C^�͇��$=r�Ҋ�8ïKvCr���{�c�>oɔX���n�U]�ý;+�m@J�5k,D�N>uylJM�O�칹a��,omÑm�����Ny��J��K����y���`�`�.�埽\D�+t1��A�Et���rp%?��l��Eb��/�n���tT2�-���`5�^A��S)'��V�"�)�;�h,�İ/��6N �7.�,!��,n���GF�)�&��>��W��t����';�A~�}��o�Q�ƽ��3����D0�W.�ADBr� Q��r��aQßƳA�J_���`D�Bۙ��ჲ ?ηo��%�3'�?	%%G9��q���=�Hăf�#Tߺ068b�[I��n�#��	�\�D'.�9X$��cݸG�p�����(:vsʞ���y!�*m,:���z�=�A�V�f�FR(i�q��o�t�6������,����PU�֗�ϐ@A<~~�S=&`9?��_���^Qn"p���h-RD͑A�����Y��c�4�kק���oA��;��E��f|q�0�i�!���6����?�h�I�Kе����[���6��X�6���%g�r�Pv��j�^B���C����@�R��B[+N����3�n��J� �:�%��ӭ���oor������B�c�Rs���0N�V*� k��^�za��v����D�t�>��	�9N�,`���K� �&�$���5G��hH�#���'K��2�����@��3+P�p���y�e����(v,��o�_���¾���r+��/��X1W�#j��j�>��k�-Q��)��1�N�y�aA_���:�m�>���׭(b�B�E�ܰs�9����W���n�=���n�V�lg��!��yeq0�����hrZs���_b��ba-�guJ�wF�Pq��W�r`Ǫ�FB�(��������<��g���� ���dU$����c������u��;��u��JR��M�w�fCA�]�2�B:hӼ��V���g�N��2C!�S6��R��rz�݇�6/��L��s^�
T:�t��q�TC�/����4�8�ɷ�#	�{ycY�L�ܴʵ���B�o%=�x����y�a�_�gVz�	{��Jq�&��76%Au��Γe�f��*y��+J����ޛ�C�v��/�R��"k�v$!�v�J��mT��'�蝢��(E��}�d�:�Pc�f�f,�;�K����������������s�s��s�s��^���_���J�����I��ƴ�:z�U����7�����q���!m0D��ݮ�蒖��c�m+����-��7+��1�+u[/R"���7?J��9����������r�L7YU���iV3��(9
{���eK4	ӑ;�j[�@���gÖ��}����Ӛ�E�]j����Ұ���<�-<��w�p'�$���	���cac#c���x)ϣv5+�O]jf�X4N;0�8���29�۲���ڰᤥ�y�,%�S7<��M�xX6��s�1ګ|������I��שּ������W�����ː�&��r�]#^FIjGc���s
����uι��׿�Ե���Xf�����s�d4wE��g����U���1�����~�~�yc�9�W���skKNn���2c�pu%�c1�N�HA��s?o��c��3�*�m�z�ޕd�3�,��#�n���>��[��[��b8?z��3�ĉ\w������_l�.f<O�g���B�/|���M��۩���췍������ٺD�ܗ!	�{j� �ӫ6�Q�NML�9�_�Wr�*�f�is�I�����]��D�U[qf2h7��c�"���@��J:>yCx�`����9�/����.�w��pS`�>�G����`b�C'6�W���;�^�E�Z-VY̭�w��JF	=���9��\�`�]���'��5έZ�~A�����_�T�|��o���˿�[9��f��+�T.�M�y�^���%�mj:�����cOC=*�<4hǚ3���b�K������������ ��g�W?�ѬΝZZ��(�)����"�o�-K�W_G���b�鷞�O-�>%��n_O.��y��.�ѝ5}=+u�y^�/s;�d���˸ysv�Ȝ�7G�G�W���S/�d
b�����oR|��Zj�m��9���+��:|�Q:-7����_H�-lq��~]�ċ�W�_y$e�L�ڜ�Q\�Fx�=J}z�zۅ��� c��Su'
5����7_�q/������>/�� �
�L~�O��V|/��I�umEՎq�1Z���|;kM/Znuk_ؘ��R���Tt��|���<a/LF=g�����0ۻw^�1��>���mҾMR;�ʙ���q�C��Y�22�a�̤ꋓ2����Եl�]U�X���=Mʜ�EnSq-%�Ѷ���%�_�yP��~p�h-�zF���
�Lb��N��	|�n��^�l×xb_�I��;���خGR��_;��m�2կ�%,f�i���{����ޭ��n�������օ6��cY��2L&J��!�}���i<8T�M�΋<ZDiu�$�Jo�k�)`�._����ܥ;l�n�OK[��)�O7��X�g�����D�c%
��Ԕ�{
Wg���UZ�՞�zc���W#{�9�ch�������?��s��L�֙z����C�����<�ff��u~������|�$Ffc �hڴ/�u����P�z�&֟�m(���)��9ɛ�ǧ�Ǉ�J7*S�+ޅ݋�h�­��g���Ͻ�e{�BOY:^�%�D�4Pƽ��N��}�1_��r޴�X����E���*�u�D���&_,�w%s2F�G�:�:�ޏ�V�H�+髟�[5��>|e���dw�Aj��)�8�[�|�O����~�����,+~�7Q$���/0�
Ͷvb0Z�F��cV�ݯ������ӭ�~��Ԉ?�on��B}��i�d\�r�s�q�}�E%�i����4��Gj����W]���[Bw�����b����D8�a!��5�v��w�V�#��hˀ���}:.Ǘ���Ɔ^U���4�J�}˽�.��)�y\�@�\����p�(F�1ổό�ֿ�e>V>0����4��묤�y��d������O�υ�=
�>q���zR�5��nP��zV��۝h7���S	�}�KD�)�ǧN��#.\4DT������;�m���|[�@�O��f�ǋ
�{S������?�A��xr�u�I���~��Ĩ8�����p�۾�z��и�b�X��l-|�}T�Jyf�\�(��[�"v�R�vD>�~I�H���x�k�<�$�PT�kB{\M���B�]�N{�9]5oiRR���YY?�a>^#���QL^�N�'M[�E]���:�:�g�����6^oZ�r�y�'b��aY��s�.�X4�,}���ihbK��w��y+��n|�>ʵe#�ofO���&�a��ΰ{��>h �L�>�>	E�w���n�9���6{�
�o�3�x�L.��wv����7GDb�]�z�a��n�h��3-���΄x���.�/�ʳ��jVa[X�.�<�,&�q�	����M�s�{���s�aq��a���}Q�O*6	��n`���T�d��5 ���WeW�
�	�<��{�����ۻ���g��Q�y��p�������[��[��7�3�G�_��Q�*��;�P��_���z�s��g�C��E)Z�Q�o8�J��eS~�Z1��o�Ck��n�NML�ۅ��v��]�d�_y;��6�SnI�A��7J��K�Cj��1��sԖ�|.��Yb�y5�"߃��__�ל������O��Ӊ�R�#�E��Ϋ�ʧ�������i�ī��e܎7�b��Mc�h�����myg�6�7��hR�D�,l�^�����S�l"��j�_�ϳ+����&xwj�g�v����ô?am(�`��	�]�񦀐�}������ߺ݇
]�M�����ɠ�h���g��O�8��+�?s�z�ݪ��9�ߪE\��w)��9c�7�0��ϟP	�O_�i��ƣK$o'^xh�S���P�zN֮�|o��.̒ߥxw��y�\�%d�i�H��/و��G����g�6?6�b�.SYO'����wj����+r���=�<�홱�K�-�Q�O���s8Ɍ����Q�cKʳ`�Nx$�g����������U��#c6�������ʡ[����v�K{L��)��Mt=���܆����$���ك0Ҫ�����j�ɟ\�;+s�b�SG/
�,��mU���V`Wf�������>_�x���iv�.���_{�V��Hm�K>����j�qS�����+冋�4t��t+�Ժed:�w��hy!g�'l��JÎ��.v|���wb�/N��11�q֊����=�Q�6��o�vM������ҷ{������&q��^q�iDA�8a^��>�������և�*W���I�T��k袘��Ч�,l������Rڷ9����i�&����wO�ND}r�{>g�9z�i���b��D|Xe��J�7�=:��/jlx��!y�x���r���=�7�YR����/(�������������\��ϧ'�vPW�����=ee�t�x����i�~�-&��&��(��/�p������ZZ���9���a؋�k�Ԣ��͙뿽��4/��h,��\������'���VR�Q{/��Z�IJ��Ms��;.��^�)ǋ�>���c����g��]5�ʯ��L�c�U�>�j��iv<P)��_;QW�n�?�պ��n���%G�I׾���r�iK i�����}/VR���C%�:s/����x��1g	������ôiK�h�/�����oJ����)�X�9:u�{u-v��pF�s�{Ea�7Ocٚ�9>��M������]y�8a0��#L�hʱ�o����NOQ'o��.�����S�z&P�~�2]���l}��F>��,��:��S�W�7�U���u�V�@{!l������_6C�+z��<�V�UⰧVR���h��ܫJ�B��ˏ4�q���|0�m�aȾ�ݦY�Ǆ��)��~sNȸk�(s�Yu���+���z,�]���|8m5K{�H��Z+j<C��9���n���{<M�X��>���Ǭ�W?)in��]���&�w�'G�e��äx���;�rb���!;�,�{=l����}�@�\�IW7�}��㇬�����F�����SҿL?�n�5uַG���uu]mZb��.M�9��T�zj�f'9�^4����B���P�/��x�����I���n�@ �Ǒ N�2�3iM�]}��l�UM�*q�Bڇ��ENF�:�{��o[�-m�j�j�~D��l�fzJ ��鋧~�+Z"���wv����w��j�7�#� :�~�a�Ah��i����D�+n^��Cw�Y֩�����u���xmh��[�D�o_�ft��H����J��P�X�D���!�~;����Ry��{����M���ڔ����'��G<�Y%�?nlZsm�Z�'�\�j���{�Тڏg��Ҏ���W�?nM��ˇ���yn��6U�vEF�B����^���T��?*�>ǣ�&Ls��D��ģ��'��`j2���g�j-N��u�z�\^l��+�0Jk�����n���k&���7����T>/����k�e�m,k��*�a\�^�w�~��yo�%�Fn�K��{��e�<N�%��O�V4��n?�\e�d����P�=��6i�>��,ǔ���#���~>��{�ޕS�#�G�G�)sJiM�m�վ�����ΩՁ�Z7�Y]i|?��v���}oXaY�9y��O���u�7�m%"9�G�����<��ϧ�N+��t�MN,ʌ������_��#n<��l��N1�l�ٱ=p��*OK.�8I�y�$U#��N�<�ױf�i��*��oy\�5M�s	�~<]�){\�t�S�C5�uO�U����㭀���C�yJ���������A�+�ۄ��=,�_�r8e�v����q��Z��o�y��V���r$wqװ�j�q�'��,�\T�I��\X�l�|Fv���ւ�L��.���z�Zb�r�Q
ơ�g�m��nX���9�r����m�����+�]
U�t��xS!�v���y�g5/*��ٟI��yɹ�|܇zi,+�'V��q�}�e�Pv��f,����,��`�Sj�m����;>7�~c���MYⷹM��~�(��z�������s����S��j{P`e�ʛ��)G���0��=\I����"~3�n<b݌�3�L�tL�*	��T��������z��\]W�<�(�����^�������?�:���xH�P�u�T�V�*�oK6��T`#u���̭�:�m���h�]9�X�aE:/q��F�grL-��4яK����'X~�����䕯�+$j�~�<PV`S�z�巀߀�E��N�\�a�g{&I�_�ϻWǗxui�L��g��Jq0S����l�!*+<9D�UK#�B:pz�����}�v�ҿ�<�:�3�c����"��e��p������_Yx���XK߮�����g��iK�?����Z1<��[uQz����Α�ŏ�kK��iO/W���ݷhI��v��gf+7�T�d@��	�~��4oQp�e����E�n��Gm�U�X��Y������d=m���✞�V"�QV���νg]@X���Uz��Zr�)[��)�ȁ�h�f�C��.-�m߼8Y�k΃K_%�ww�"�'�~�p�d��C"�b��зCw����*��/b���w�Y6�����V�S�g�X�0�حԾ�*w�����W��H<U�#��wa�;C�`����s9�F_C��za�����n�O�}�p�V.�Ӕ(�T�YwC�?1�E��oV���9��+Q��48LZ0q�	��֓�U���#�G]w����*�׾G&X"���󔉏Q�0h�Y��S8�A:����TT�ٷ��<x���C�o�o=�}��C5�SQ��9P��=	��*_�<;r���˸�����j�+àw>��+�vh�?V��Sn�>���<�\0��9����u��EI��}=^�=�cѣ��︝y�?٢|��`���w%lҤ��N�����,�A
۵$n�݌��94�-qx�S5�p�BՂ�\��&���W�`�Ȗ�m\���zk�M��O����}�D���o���Q\wZ#�];'��8��p������V0�z��{U�Ò���
F<Vڻ��m�݋_*'2߯#�1WB	�%_䵙��׾DX��>vŻ%w����q.�J�Ej<6@��y㺮*˛~���^�#�x��-凛�{�3Ft�ɒ]�^.�崙V�e�IR:Ń�Ld�:<�j�ߦ��r�U7�!�պ�J�asS�q��7��?�xb���Dq������o?����݂�'ory��܊�6r�I�%k4ɍ�D�x�MA~��������_a��d���ݝ9��5�򫬞��c�����t��^�Ԏy۵�ڪ�:���H�Մzm����5]r�C�X����|]X����;<��>+������ɟ�*����Z��Y@kJP?2x����Y��2�����,J:�� �:��?�t`*-��Ӕl]�azG�`[��K�&M���t��X����O��͡��ބ��=J��_rM���FUKb�N-���?�T�`?YW���)p1Xb�?c�ܟ3,���g������W�NW�j�M��'�.^f*(�w^�?���XU���k~�)�o-�ǎ��1,O��1�ʛ"�b���c2�Q:[r�{�h��_�"+�}Mјؘq&Mc��-�a�kQ��N�[���bsE*��o'������|֦�=Uje��S��8�����his����֕�W*J�
�jj�z�~��d�%t�6���EG7`�<���&�.��bYLx2g�{ұ]�:��/������7)P~25�Y��u�����I�������;�gH�z4���"~�s���?�jv>��#��G���n4m�xt��������\�+ϥ�9O�~�kH��>��ٴ���O�5��怟Ϲ�Jκ�C��E�(o��mO�p�b����V�<q����?�����F�%��.�U{6�-j��{�r�M��VEo��{���-k�)ɿ<����[>s��T����x}x��B�BE��&����oW����\-���l�C�j�{�0�],{Q�&���%\�Z	�d�Hϕ6�n'�難�MJ��!R�/ރj\ZgI���.�s����s�m#+�O��7~�i9��c���h�/�d�E�CԆ�^D���N��i�ɋ��8�~��7����\W���7�\��b<�Xy��
N�v����מ3�A�u>�Z�ɣ
�����)0��,=h/ꜻ㜤�ܛ��~��-���:H�a���1�[L9��;����pFzK�c�=���J~S'��q��b\�M>Ƿi_i��&��^���R��� �*��yi��F��Ãu��i#6�Y�����l�=�frTQ��;�\�!x�/`��'�؉;?�o����F2��W�f���d}߅�;���&u�|J��RL��'�|���N�k�kT�H��5V�B��o���{b���k�+� ]Wqo._q�<�ڻ��Zb�O^72��S�-B�^h��3aRV�|u����ʊAOxP��S�4y��b�L�"�l����e��#�w�f�O��xq����hJ���I��}�o���]�� 	�D?���s�;�OZ<L�~�W����+�A�ІҪ���v\[���=��4�Kw�i\>Ns�o��yi�k.@ӺO��0�F��=�t�E���Bs��q��OMmi:Z/�ۥ��g��k��S�_L4�|�L^��k<�"��r0�͡����$�P����H�.��&����x����J��-YS�}�m�5.U�K�	Y2�D���K���/�W<�������o��
��{gB|�$I<�?Ё�S�3��[����Q�ɱ<����]�k!�1s�c׮)�u��x|&���&�u�V��s3�&6��L�5�q���#�f�ՉG;"�]�w�T���M�q٘�>�w�H��k���]wr����CVO�>~>����.��K{�2��X�����N�>��n{Ɔ����r�Ǹ{z�a�4:���*	���)��&��&��Ð������h���Ӌ����R����oL��?����1-WC��rW`�O�Fs-��7׾�<�H����r���8�|N6��vO[ p
(䍄�K�pD�*��;�n���\������3�vefO��n*�����蚉$�49v�t�d�c���Ѻ����[��������<xpN7�X�/V���[(C#T��ڏ�n���L��е��Ѱ�\!�R�B瘽v�l�&�����w�Z1���Jo����菻����%��_�'E��S��	����[��(�*�V��5g�IP���y��&/��W��)�n;���e�o����m�"5_$T_K�?�k��wd�½w�^��;v�����.<Z��Y����M�+��l&q��K?a{7�kR��:����Y��1�I�B��W�_�헒W����Lm;3�>f��n���wK}���KJl���Y���)[��OM���s�2����ύ9%p�����s1�s�0+WVVn��e#V��8�K�Ju�Q�}뽂�jw.[,��>�l�΋!�:&����ȏ��fq�CAwf5?�$��شcC�≟��޶`o'�:��6�����P��/���h,&�Z �5��K�h���xʌ�]�񂥼��o��<{*���JF�A���鈸3R��0���0F9��fDzi����T��1mo�,E�*�B����b�^Y�n��D����{�`�8��'��cq�R�)9!�ܴ��/���T,�����Qj����q�z��1J:���ȋ�M��Kz�J��MZF�b����J-5�?�M�3#E�1��<������SW���ˬ��W�Ͻ:\5�9�����k�W�t���f���kxTv}Kh
���1��������1�|sB�U��I	�ʋ[�4e��܍����ȍ������,��ӵ�J����X��0 �Pvq��阃���ƈ["zx���s��n�\�y�']u���P��I�q��;����L�(����ٙNK�C;צ�S���\*�x��ZX�����R����������$N�+���M9�k=���x�'�w3Ft
���Y�Z�ex���:�E��F3o7Dϵ�0�Aܥ�����I�z��_?��1ʞ����.�+��.⣅.�)�N�n+#.n�k�,�@㾯�όj��PFTdh��0������e���u�bo�3ք���u�1b�GtX�i��e!ACؠkP��H8k���� 
y}xb]����`���,��fj4���=u ~�#
�O���X^�P�d�F�.8_�{u�Y�������~��t��"�#SA��IvF����X�kӛ�����v�e���<�j�ؖ�(���1�4?�����Ώ}L�"�-��M�<�zW@67'n�}c»����)=��*iکup�x�:')�)�I��3Η�J�	���a���%*-#�5|u����K���
�,�.�Fë���;�0킮o5n�c������|d���=˓t�!��?��|4=��d5T�n�ƺ��V���5oL�FFds��fh,t�Do�_`�;Kk~�2zk��,�s���H���&o���u�Ē���Z��0'4|^�)H#%-܊wBesٳgy; � CA{���i�&�[�b��@�'��s���כ��|��=���ҏ�<e� V�ЧI���;���ٟ���t�3��$��J����l��n��j�0+��^ʈQ�>�2t+��$�J�#��CW��s_�� ��D!_����=J��Ҁܺ�+4�Fޙ��@�J0$ѫI_�)8�X[#���Ǩ��}1 }��d�p#�h�ff��s�}��I�*$��e�c�SO%7m�����l01N2A������涊m�sb�aa�D$����ey�?�4yH���N���?{�0�rDo��I0�m�vo�Լ�*���(���g��Q�#��W���܇�z�]�4��M��
�@|]��1�O�����ِ�جB�;0��L����HK�8k4�a6dh�� ��Ak�� |������ȳF�T�'�����Sv�����ќ�h*��]��Dl�m X��/	����k�1�ȁ�Fx���#�ťqi��q8C�hߧƤ\��^}*|q��D!#�?߇r�ء�ɇ�Ih5�۫��uS���т�U����az�BQ5T��S�6��o&!���?��x���>�9彣�Y]@>:��1iD*��Ԇ*;B� ^��E@o����s��t@+���=Ϫy�c�V�mձ
�a�ֆ���lH&nw�sr"GtΜ�����0�fD�q���X��vd@AJ�s���Bt��S�mD��[��*}O����e^����~d�� ��@|"bEY)��Wֻ����YnS*����|`1e���|r��z�6R���lj�W���8�Z��~���������X�s�<�{��:�p'����Ǆ|9�5�8�(�R��hG��?�^>�n�K@��{���G��� ~�T��+��)`�"Gr.�aj{�Ėd�i?}YiF4��:�}�ⶣ��!�[�f�}o�P(j�[oޜl��P(�P�3z�=�`ɢ	r2�]3��s�#Q1����\wv'JR��l{� f�Y	���b��/��O���wļ��j-�߳�l���٪3�@h�V��!�#橭V�>�Ě�}����=��6�Iy��ȉLZT�b�w�	A�ڣ��Î�x�IpP{,.�(����v&�=|8�-����X��J5=�퉡��6�n>�����5�ak��ຄFF��ng�=�����Mǭ�'��O%��)`��ec��|V��#�'I�b/�x��񷿞�'���D�"L��{{�'����lD�3����S�<vsߍ*�j��ԓu���(��ܩz��+U�C�?��P����폸u��G�޳]�JBv��H=8.����}�����S�A��9l>�D�<�w\-�t�#K���������"#��S\G��Z���=�u�d�r~lpI�����G�aO{��ͽ O���B	c���@��o�a�d�#��j��3f����}tƿ>vcVaVaVaVaVaVaVaVaVaVaVaVaVaVaVaV��z�?
����/V��V�.ۯ"1�A���^�;, ��w��k���:�ή���:�ή���:�ή���:�ή���:�ή�+Zw6D��(��t�|��~�vv�]g��uv�]g��uv�]�/\n���׻ �_�2�ή���:�ή���:�ή��6g^����\P�g�gbE�3驖I�Yh�&��-iJ�W�������*�MƼFtc�=v?�u��k����_���j}�bh����z�Mm|����l�g��+��mg��50k`����Y�f��50k`����Y��_P&ߘ��d���7���|K�<��-���(/'��v7���2:������wb�wI���|/����r�yc�
s0ڈ����	O�w:�������ʊɦ|^orDor���?���B���RxE|�]�,9�:1y���C�)F��0�ɸ��?��/��,��9o�FM��:i����i���~T��b�\#�{OﱱŒ%�e��'*����0�'>\ՈY)G=��-�H�X���I�*�������3T�W�| _��WQ�ĤFA��x�~�DRY����NL����jIc�b�Z؇�T���Pu�z�&����X��HN�b��е̠"dF�,*��r	>�� T�w���pib9��nvb��ɸ�_Ȱ2�����&����߅?oUC�,E�0����y��|�퉊
�󏼃%��Ɵ>��iQ�rE_��(h�ہ}����)�7���|P�F���`&Lp�rl6t�P;'I(���=�`�E%��~�O�����{)�X�](_�F��f���N�r��\��kޝ;1y'׼���2J�؜��ڠF�ܪ���&�a�np1�/ӡ�1"�
�n���'�Q��Ȱ�,M��l���Tx�(�����%��>���?�SL�u�eQ=g,�∽���qΑ��Q.��!���TB����.��$����'S��R@ċ�	�G�$� e�B��(���Xi��sl��w�nF HB��y3ԑY6�}9��t�O����g��%N�* Ჷ�s��n��#��+�3�#_~���>�3 F�#n�Cʼ��<�����]�[�!�`�𶙡0����%`�O�y�ϟ�d(#�5�9|r�)�3S�?��Kt�Iq���nHQ�*��ݽ	�������8TN37�D�!t�7����l���q��p��~Ri�yG9��Cԝ�I��2'�*(�Q������F�, "r��Vt^)�/���-�����QVe�ڂ���D��%ePbMr�T�2�&
/���$�d�Ex5�����L5z�ո�����Y���Ah���f(��iAI�1�t��oj�ā����/�d��#da�'Ya9C���`)�K'�Ā�5�#�QR�/��30
���L��ڸ��tP ��Ӝ�IBT(��)(���q��t\���ÖL�I����� D?�J5�K'�.�U>1�d��Qo\�+(�DdREPܷ�<Ce��U����� e�T�V� �ԮAҍ֙��.�+C�T���Du�#���w��2��əR�t�֔���݊	zc"lT�:�����b2Ȭ�����>��C��6�s��U �Np3�u�L���Qg')�ŏs����nO�Q ,�`41�H�5� "�5�Te�L���	FʕO'&?ч�>�\+} ���F�L-��"����F�́�-�ٱA�]��WPg�D�VC������98�﬎�B�Q����3G�w�,)Q;<4�ϟ��������IK�0lx�>s�l���������N��V&��57���!��&(7��L��upX�ߐ��d����q� ��>SC�zh��w�ߊ�0�3�^�A㜭35i��12��*]?�,7�����wa�S� q�Iy�3A�v^E�P�2m�;ᝉ3ѐ�
L��͠�z�D1p�DA_Tğ�NVf�Pј��)���qj?�r+���(Cqa?�\�.=�u�M8Ȕ����	���<�F?�PCE��qxp�L+�Mx���H�S*d$�q��������d�<.�a������o\
�#�`ɝ���qѡt����X3tdt�#�6@GF�؄7�#>�
N��J��������ѱ	�0i�DV��Б�R�<�����	�+�^�A;�� :��������ꭔ�V���̡k��Z�2����׆f�<8�C�����:�Q��@����q���KG�A�Aߔ=�L�+��S
�����F��[��鈎�@��}))�a������l�����«7�5���u�'�53t����Eo��a��T*}�����I�����|Vv;x�`�8������h�S�+g~P��4t�I-U��wH#g��ۣTj];Q��\D�}x9�H0��; mF[d���[r��	� �g� �� �_��'����n��4���.�1���H#_[Qa�1��G�Ժ���]zR!�E���O��U����Ol�~�K%B� �Q�����2�5h��-e	[�bOQ�����|�O��>�Z�'BI)·r8n�ՙe��4�_6T��Q���&�9�}����� ��^8&o�N3�������'P����g\���`hC%�}��%P�i3���@Q�l�5�m@ABܘ�����م�l�ɏT��Yd�@����cXLPv�#��CVW�2����d�eP��N�����f��pP�gtȍ�ƕ�����������"��YܸG?��ɹ��?C�S!��wg����J�C��-�h�5�!��yS*���U���ȡ�D����C>�T&���^- �&�V�7���'Ɠ����H	���ߐ�^�E>5¬5�v|�BD	Qb$n������/�|�Ռ��F�r�u'����\���F�y���7/����F�\�An�z����qo|*���$���+�9���������36;�ȫ���p�re_���:~R��D_������v�Ers*g�s����G�f��L�N�HS�D���wKQ�%�@���Ar`���ޕ��Gy�����r.�.B%��3ݐ��?�a?@�o�HmӝI%�t��oVָG��S��:@u���%�� �����$�c&MG����Q������g�~�x��b��"u����
 �9�34�T�r	�����3I߹&��1��b{��w�@��T�u�f��c��ȑ WVQ��19�}���)���:�|~/��;�zO,p�#����b$��޻�=`���zo�z������`��*��,���\4�^9�Q�G��Y�ȋ��1ȡ7�c�ģ�NTQ��,�s'�5h�(TU/�@(��J�	0灛{�I'~��M0|&+y�����>�N���O� ��0��Kj~W��$a�'�L�K;QY.���Uǰt�O �*��~ �W���Z��_3�F��@�x� Jsа8���%�Tu A�Y���p�ͽ�d�!���2Q6�}��d!��O�42@X"��M턽J ��d���s_S�׊��A(�(.�*�^&C6CR,�2l	#MG(]�@2_$�F�ޢA�Yr�0���.i� 4<��R�W�$�E�!+]ڎD_A�;�u��Y��h;��N2��:��]����J��!K����-c���"�!��%%�ˬ�;�ډ�o�{õG3$;2(�U�b?��$F�#�E*]r��fGجQ������߲�BBpݡ�f�:K�&� slD}3W�N�z+~�D~H����K��sI	��^���.)��ώNm�{��=��܈z����F!�A+�Cw*���fT^�p�3�	z%~|�	y���M�#ݸ�tIl+��c�� s����(�q����-�� �����qX'p�n�鉁��>�I؋d�H���2�e3���Jګ{=X-�[zs��Q���Y{AF�A�*�1��L؋���n{�,��{�\��ڤR/s=�HF2M$�YiSK6��#���{7�#{����"�˼{Af����D����Z���)G�"^����\�'��?��"������b��(�%��rȗA	!�B���U��2�f������-FSR3�w��@0#u&��9��߼�$6z��KfX
��RtĎu�&"�:��f�����tC��9�̇�v�._���X	-Qף;@�r'w�є�:Rż�Ԥ��"�	|9V(ƕ�(@��^��IG�a����8���蠨��h�$�1m!����=�����A,�B"D��Y,�l��� �1��/!�_���5��)���|��Y(ʖ����I�e������)�/q���;m���QO2�iY^�EV���r醌�`�����dt�T4���yg?�_��9�~��~k۝Qhs�P��Y�12Y�2w����b�e�a81;�)R�@syM�q0����G"� t�����5�B�`��cq�d3:j/�ƚj?B>4�e��C(��HbO�RC�E$��˭�' v��-*4,��"�hX�Pǰ�)u!��Fj�j;r��5h��f�Є�(C;Cmr���iY~oL0h�\I�����a=8}M�VDZ��Nk;�p�7�S���BC��Z������s�[�B�nPAִ��Kj�3=/���N��9��(�Ks �	���0I,�-u�Hڔ"��8@j������1@�����~b�0��Ajw�!���?>�f� ;��\N�I��H��U&��&�r���ć�*b�~�Xp���A8P����zp� ^,��	�p»Cd��^��l�����^���_��K��[�����(�}/�H#��؉~œ���!�~^*�sA��S��,h��\W"��,-��q�A}��Wd�w7��a3�ڋ׼$W��ari���� �]�"]��L���D��כX{H)��:N�"�.�T�;,sp
�&�#}j��R�Mkp���a/��Z�S�	8�pk�AMw
HW�2G�i8ő�5@J��"�ӹ�S@*����zrZ��7t�HqeM�c�^й(����C��q-CK�h��ʐ��A�l
~[��&4�cI��V�HQ2��6��؂�]d�w�.�V�܏��7�2ut�?��&n�e0���2�g|�B2%\c�[-#�B�3���yK���c���{�'��)�Ռ>؋dx�wܪ������\�^�7�} z�^3<��2�g~�B2�P�!e& W�h���$;���>f�}z�p=�!B�W`/��ؚa�2�fx�^Hw�M�w��e��^8Z*O�L�5��=��C�$��8��[K�z����G��K���83c_�l,A� �%���6���"��4���1hkt�}�YZ*�*��V�F,��%\Y�}�PH.idN&ƪj��&Q���Z>���A���~[ɕEe���s�K�, �����$�md�Ҙ�AÑ��Mn�NɅ�N�#�c��M��c������O����K"�2n�\ko2�[@�����������<#�!	�w��&A���B��&h�� ������jЂ�W��(m���DH!���@�f��3\�fn�� ��e˸�P'�=^� �N�8IL'�j{�n���B�A(�^�s��'!��pԗx���9u���{F��qV��X�c_���I�J��C,p����]�2��B%�b%Jˉ��:�-�F��������z���<Y繲Rz���	���1(R�~��bh�3zWAoٍ~0\���bYxy�37G@�&�b�߁�*
��r���pG�.�sWֳ�����y?��k�O�E��`?�w���rsą���%�2D�I�X
QO���|�C}���M5s*ʅ˭u0�|-�:�0R���ڶ:!�C}%I�R��\��-�6�ؑ^�+��g�Ok3K���:�D�#�B3��Ϲw�Y���y� �t���[��[qcB$��>f��������^�'ޮOQ_��<Q�80�E�o��Zd�+�<�́1�Hx®#�����a	0�+��a>ai-��E�p���a^�e��~^�m��0{ �2R���f��L�$���90!�Wq�4�V�K*��i�8�S���B�r��0�?�������p��'s:��ӾB�T%吡VѨ�-Λ�SH���:$��>�"�
�>������,�H"p�2��V�3��(R�/�G,����A2�~�xH�w����J�*��'���~��$����%��`j�^����
IR��]���� Yx�O`8d0�,��Ӛ���u��Fh8����\�k���[���Dϣ��W����-�㋨[�}�+Ε=_���D&Ae�!��	�P<!�'!<<�����܈��U{�m%����֒�� d8�_����|(��3�6E��[�Z;�3�Ǡ��!�>g8�{�nPc�!��N�A�((E)�f��j�sGw��!T�<<H�Kkĉ^uB��7�-u� ��Kg}QvE��f���X|�s�(�-<���_ο�w��";(�Γ:���҂���M��e~�/�
��{������J�Q���:g�l�5h-P��xi輦~��F��f���,��#^����rYZ^��يF�<nP�+;N�E�\��"���@��A��=UÀ�[e��F�z�3�B�mB 4�`@�g�A�N|C�*���ĩ8��,-s��-�K��{��b���rnD4%�4��@0��|�^��ږ(��
-nY�,�3q��XZ�H��e~ځ��f!W�g-#�>
�p=5�{E���-�ӎ�e�Ұ��~��g\O��'9� �����_-|/t�F���[8�p�p��,������O�$�U�����ވ��0x8�F�t���ކ��^gY���kv��/�!��B�����Ӗ�v�[H��Ar�vnD�h�!E���E�#B�=K+E��y����zrT����<�^g�ۜ��M� �G�F#���FYێ����Hb!}Ή]ڡ��tfs�3��K����D�Q��J�ڐ��(,�@JG_9�r��"r6j������@�1�"� ����#ކA�)�PGצٲ�e$���XQ��+��b�E��r[�sO��9��>�=�yϹ�f�n��R���:f���g�A8�3����Ƨw���s#$3B�N�_���Ƭҹ+�O�W���@<��� �2�* &�u���UR�w˅��Ư��B��)"�I?%��g��{͊��y�sʂy�CB׬�OȲv�ID��c�aD�����R�O\Ԥb���W�6�����S�^���g�z�=���E�B�7�j���a^�R���0p���M�WlQV��*�K�?o�>��{��^�g�
Y�Z?����9g��Ա ����-ɏLH1��A�WZ]n�M�8�=�]��0h��Xh\��
��3|D@n�o���u)�jd�i�������R�O�!��t����Ъc!j���'�-�x�ʜ?z�ڏ�46;��|<�������p��;tE��p���t���f�_����nu̖���+��u�ަ�cs����z���9���T�0�V����<g;b��V[Ƹ|Y��6�a��QY�$��x Qev-m4�h�,�@�q����S7!5��g-�7�h���̸���dÌ�cxo���`��|�]K�R����º��g�
l��3<�+�Sf2+bhU�Q�4�zݤ��+�_��u��Z���R�a\1H�����"RC��~	�R����ٰ\������^O�&$+n� �Ld�b\�,\ i��)5�J_����ŤtJM����f����P�{�\o�R2t#�e��ܪӆ��\y�a��];9��g�PK   ��X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ��{X`�/��1  �P  /   images/e80f2fa1-d37d-41df-8a09-120fd0c34151.png�zwT����ke�ā�AADz���F�P�B��5�Q�T�P"��@@�@t�^BK"Aj !-�=�o�[��w�u��ho8����9g?ϳ�w����/��� h���!h�$my��V���vI�����KA4�*����8>T
�s����C�U(44T���~A�?ܸ��Der-�!ht��{簬F��١�+��
�폌�TtXjC����ѷ������o���n�щ}��M�^x�}�uWͶ�ߔ��f�Ǵ�;n�~�Q��W��z�4���xŏ�C������W^�MZEǰ�1�{^��9���Yne[7�A� &��{.���u��}[bwI=�"�<n�l�lܨv��~�i#A77o6���ɆL�1����'MR�%j�&����!�4�UF�u���a��U�(��HNU/�"4���`G��dN������z��7T���9��\Č�ق�=eOu�Z	���Rl�ƚlGXYQ)��oVu����k"qz�g9P�4��x�T�ͳ�5!�U��i����#�-s�.�	�n�#�o�P$|Ek웅ĊKoE���K�-;᫞��H���f���0V^Ϟ
���J~��d�5ۙH�^��Qɿ=�Ƕ�%��V�._�|ǽ*?ͩl���-$n)����.mY�3���j�q�0�6��Ŭ儁��HSH$����m�ȥ�Tխ�'9��U���`�J�G���
w�(S/E�4��j��,�/��ˠl�����1��P//+n@�:�TБjgP1y�q�A�m�Zhs�03S��k~ק���SM����~���)ű��ٕi�A�rr������a��Vi�Y�v�iy-L�KTD0��B ,a<g��~oBnr���`[�R�2|�vQ�%��[��f��x�ӳ�/�D]q���;3�P����̿����b���0�jy>i�N����OX%���D��5�Բ���F���SI;s��Mv�qV��.mۘ�/"�,'��ʸ�\h�.C]�����i�ײ�ͼ�P�x�|FeS���K�f��(
� T#'9��(ٚ#uΈ^M��C6��c�?��1�4b���?/��V�*�c�h����x9�Hˈ2�l�1:f�C��ժ	t.�`���8'rVs��ޱ-x�%�X�_��ZA��>x���5i��©LU�
�{}��X|�H�뾒,���%�U�K���s(�������2}����:Z�+
����*s��,
���Yl�$��F�~۹	�2��	v^׮�s�ά���;5���&�0�+"ѥ+rm�ӑ��1�^J$i��1g��1�n���i=�)�T\?�V5�ęU����(��������öfo��dG�%��mmsk�KW�dii.����N���^�5�x�$���5�Hx7Eֵ��<�w	u2YxC=�~��%���F����	��e)�I��~�w�#"[�u;[g�C��z��ZL^4��Z�V��v�w�㬚{{ Q��/��5�p��_gp�0a��9����b�4S$C2^�x'��DbNg��e�w��I<���I����n�p���ˢ��hsl�W����!o��s�����)|�OѢ�t��؛�a��ţ��U��y�>�GzEN!q��\Z1L���|�O�`$�I�BɆ�������{&T����$x�*����V�dڄ5$�M��Dko�tD��)C����!�5ʘ�@aK|�ׇݓo��.�'�񓪮j�1��6|�x�F����G[C��&e�~�]�R��R�l2��};�b{Q��d<:J��Q�}3����mk�
���8���9��<���~��������o1ϊ6C�n�2g�!E>�GsD�?u�mN�|�1;8����jc֭�p�����Kn|�{�3f�<�SD�7�J�jPZI�Sќ%h�ED�M��+똢��[���,���� t| imj��".�_�iܔ������c��㪐J/��ƻ{m%,�̉Hw`n6+�G�:�NJD�t�U}B�0��Z}#ҍ���q޹y(��!H�'s�6�L
^�zc�#���^	�n�Q'���_�+��W�kƌ��cf����,\�����p��N�[�����I���Ss�?ݵN�I�o��I�I������j#ꪸ����&�m�?�y��)g���|�|?:�+���*�/���8�6�?���J4����SS��5���x�N$V�Q��q�!���s�dǒ1%�48����t���J��0Z�PfbvD�Q����M�"bմG�2R��#R^D��+刾E�Um������uA}�I��
�~�Շ��S�u0�u������!��d�n�Q���7����x�|��r�|�ST��kO�d��pf�G����c�'F��adyH+y;]�Q���$F"���o�ܟ�Y�����ck[\;3�*x�X�d��VDVQ��mz��4����A���0����> Ph#M�h�ī����t��[�pQ}���YY�H��EN�����n�p9�l�Q�t�sݦPM'fc�)@bc�R<�@9�?x-e)^
��-e�^�)մ�{���4� ]y1����"2o�@`7���xZ��R^y����olP��_@[I�W�K�y�)ZNx�����^�W�c�(�����Ʈ�'6�Rf����.�o��
�5!�e(:J���׳��VK�;��`�;0�[�x�aҊKG�V��\p���n[����1z	���z���i����/�Vqke0�J!!⮬�r���CJ2	��QNG�E�_J��l@#��^}���C�]�k[�2����6��]隙�x_��`��$�ʿ�\G$�����X�f��I������Lq�H7�>�D9A��-�G�ٺ�g��Zi㣊�� �3�[5�P'I>�ּ-�s��ӯ'$��0�ϓ���quwg�����j|=g��!��iy�bf|�m��/#��f����M��*	�c�-�=�v�_�R�\�@�+ŧӳ#���=���Zq���#{��	o)

��YK3`G%	�<��2	�6(݋���|tߦHs=��L|��N�>9e-�M�&3���4�C_��쭪
-+���rc(�^$?�Ɵ7w��l��$�T:��{�=G����Ҁ��ŝ�Hn�@·[
_w<��]���%�65פ'��oA��1�&�.E@P��#�ed�u,sǚi4G'�����oWL���}r�Ї;w6ut��R���������T�HGC�_�g�����ltԱZ\�>�tHH�Nir���tq���gE�t���~�������/�o�hfn��~VT gj�������Q��m�����������QGY�S5�z͏b��8�흧���QȂ�/r$����|�x�%7��cR:;��O�<�o����C��jb���y��N���B'?t�Ė]]Jq�R�Ħ�`��_�?���+����b��q������;[��ߚ���*�:g��[��(EB��f���dXF�iA_mT�w�ؙ�&~,�p����	^�8a���^��뿽ɥ�X��(�;�`l�-匬�O�X�H*|�������[��~�S�b0�{�g�ϸ����%3˧��wZ�U_�ѵ��df��pE�����K��e�]c��>��N�2e~�B	��,�Z��ב�2�����쮦�K0E�3���/�D2��������/�w���>ы���˾�j֮[:^�����9�~�{f��d��������A�����wj~Y6��-�jlg�[/,���覹�<ԛ�U.��V�t��W�(ڱ�
LyP�N�����H:�`W�?Om^5=Ë�P粤U�
�JŷJ��4¥�)޶TbK饇�⏌��h��ԔR@P���w������k�[oę��R�8;��+Vѣ��?VYG,Q[���ϟ?G�]�啜CU>\��͢5��S	����LϺ��U��uz;a?�Ϩ���L�Is :j���c�SzM����`xDطXJ��J���J�\"�
�
�ʋ�C�#k��FY~��v��k4�p���ƛU�¬v]w�IVV����Wf�/��������t�ʼ;���ã�-;���|	�OXg��r��9^^�d�Ou\�6О\S�=j�.ѻ���B�ط$n�9ԫ�ѝ*���B
������H�ۙ�vmrM�k?�L����[��k�}Q2����i%�����������A����L8&�Kg�f$�4��2n^�'�\]�z��q�ODw����vd�eK��t�ҵ����l����o����)��̋I9�sM�&'�$<�����F6z�.l�|V$s�2Z����u�k[��6�u��ٳ�S"C1h�����_t��A,n����Ξ�R��Wk��<�_����r�y#m��� �:��2^GHq�ձ�y��H*9-9E���:�ʚKM�VH�J\t��N�#Cflo;<ߐ�r��Z��~3�e���i�u�C�+����a�^&��@���c���4�'������nW7hx��I�*�ek�p1�y\ޣ�Zrڥ����SW9�fy�{���#l�	�a���ʍGV�Ը�m��T��jL�O��4f����w`���4���'"���S��B%׵	�j����{���J	O��:'6�|�|*���h	̧��o�c�I}�֥1��*a=�?�#�}7=5�1���f��v���h�0��1��t�_'�5��jd[�^g����N�H%W���D�U��=�=�S6A7�\@�S^��I����X�5�u��.'\�G=���x"��w��n9�|��-j����ʫOfٝ�3Q#�l�9DW��	J�lX�����'�N��7|L���K���)5*��S��蜜����$؛�ܹ6�A'�ezx���Z�m-��z-;�&G-`�A����� ��*�Ls�M�����U�cA7߸��R8�Jyl�B��Cc̺�W�r@���/���G��FKo	�<���? ��N�E��H��E!��V�XZ���<ҏ	\Y��x<j?�n�ˠ�	A1��BZر�y���ň�	Y��<�%	)i�w؉z��B@؉)�����W	5���@�*n��@m�@t��%>pu��Z+��ɐ�����Y�G��t�Z.s�5�I�Þ�/�{%�h���ex�Y���cd��w@�$&'[E��a�*H��fyT~.P��" 3��"e׷��PE��J�eI=�{t�r��'�Z8$.����!�^��Ō4a��&"��d��if/L��h���W���8��9��݂9���0�)(�r׏��?m�v�ݲ��E��_�f԰D.�g�;E�z]��w^
�u�W�'�=0M/D���%����э�v�y5Ń�p�	�'�WVW�Y�R�GF`?�SޖLXP$|�2��%ZWO���C��6����.KKyM����[S��t�];lj�rkm������K�RX�Yʪ�oR���,���Z}�'���RO�ϕ^�I���s�;���.�ai��A�LJ�)����%��[��T��QG��z�)ޗ2�>�c�.�.El�>��;T.��=IaHlfȒX�賌\J%�|�ر2?zi���t��홨��G�����s;��ǉ����d �w��R �DDKaYʨk!R�蚋nM��q�vOI��`�IE��דR�p�X�p���)�-����B �{!<�yƯ�;#�H�aEP�tU>�{�	�i=[n,�n{�0�5��4������Ŗ�8#T���;?<�Q����{P�3h`:l�񢽓ࣝ
��"���J��W|��K����O�!g�9I�^M��s�h/�|c-սz���;"Pc�ia��x‒Zk[W��wQ�fۧ��h=� ȣ��h<���lA7ԱjF5�a�O}�x��@u=��س���@�(W}ҧ�U����?선,��a܈�^��� �J85sc6���[�*�D�nw�1�wow".CMA�q�I��'O�Վ��i��Lt
����h %��M��`���o�N��c"��;� ��:1Y0q���gtw�6X��]ǖ��ɹ���e�g���\�{������+
����2��o��,���9���z3V����VB��sf'��p�L�����b[� �U�iX��u�X�ɓ�+���Q<���O�RY����<P,�>�X�Щou���_��Ck��.KY��ڠ�sM##�X����b�?��yJ	�{`E�/��w���X�D�X�����U��w�{�ck<%4�V
K�י^-E8酿�yȾI�5@Ғ��8�]���R5&
����A -%��bK\�����|�SL���Fe��Wn�c���� �{��+v�1ɝ�2�Sz�/�X���i?>sʲ*+V�/�$*rXK]t�O8vD���X�z&;�7��!���f��.�����k��,ż�lj�\;��x0f�X�+a�{�$��Bҁ �������@	*q��ɤ�t������l�~K�r9�4��*0ˁ� ���%i9�,<���p������[�1��S���^_\21�&���a+��)�y�;��]����(�'?7�R���]��&BL�N��e���K��x�����O8]^]k5V�����U2����N:���չ�yف9k��)H|l�;�H>���%�ef�`Z���9���3�����X7G�����9]ζ�J?�X*�}|&�N�)��7�bvqq@4ڍ���ݤP�����;�j�S ~�@QUUZ�&HV�*�][��u�D_y�@f0�B���'���T�'F?_H�ZX�Y�t�\8��R���u,o��U�p���t���U�cj6���ܖ���V5�1+��C߂i�.%��%����n���E�	�t�[,�s:��'�� e۪fJ�KV�&��Z1R��T�}�Դa^�r����7����҃r�:��X�R3i*��d��vRZ
[g6�Q���5���D����޽����u����6���|�ٲ�G�Q:Z��^�����eC�7Mͱ�a�K� �� ��	x����,\]�r��/�ݪ�9��e,v�����^���R,sY/E5�<lAa�f ��@�u&G�gG,��`O '���ݍ��x��b�~2I���?Q��M}��8e����'۽�J�h�������-!f���*���ˮ�bl�����(��=}�
װN�5��r��l�ky�HHb~8���
A:O.�|+�a��I~�����&��[{��B��u.�3��j��+f<�\և�Ù���έ�G|�yWu
h)I�sO��$Өw��C����;����ѡ�{c���;'����uc�5)��Vs53������\X�y�HZ@������:!�����5v;�L�I6Y�u+�9ft�̦\s��\��잘l�*�T��>�	-���B �����#�&G��>�������v�l̮xR��ǆ����K_Ձ�}+���W�U�������@�NYQ��k�j`E�WZK�1=i��q:RN)n����H�tiJ:P�zᣑ/P�y�G7����u�ER���I�N,E�Geh�/R�~��v�����P�S���h��	����*}��Q� ��I�̉���2u�ku�O�e��6�ͫ�/���I��O���{���Ԍf�ϥ��D�$y6y�G\A0������ӧ��"b<r���^��J������aAu���8H@NZ��+���� �4��Ҥ�ZM�2�K��-���:iR�n�4v@���˽�v��*���o~�0���%б'ݽ�/�[�&�o��������}19s0�+���@YSZ@�E�7��oR��Ջ9$��L�C��f
�'2������6�vxmM�vi�4�������%�H!\sŃ�.��f�M,|B�̶y��}���ie��>�{�.�|y��yـ���
�}�.)��w���������n��ݳq����P������$
�Zᦙ�HOOWR#�Ck��ټ�Pu�]܏3m-�j�9�,��\�]>�_����4���R��(�^,4G'�>15�1��p����\�n����?�y
w��O�a���rכ�G�7��-�?n�%k��-d����L�矒��w��t��y ��� /����3>\��4�����5<������r�o���+�w_sv/�/,,$�v��w�y�\�����/z}{�`���7C�A��w��őQ��R�B����O�U5.�*m��L��N\$M}j��i5�� �k׮�GԖi<�%b?�^�����.��'LMM�Q`ʣ_��˫��K[F�yuȃ�ѡ~����1/iSK��>}�Ժ�;<Mxu�c{;-NNk��#wi���� IÏ�*���T

¶+V�������g�AѬ��N9�F�8:������դ?��&�:l�mh����k,SX�ۧ/���iɽ��7�`��r�jK�̥d;�%v�_ĩ�Pa|�?sͅRр��PTJ��:t֏�@��嵐���$z���RU)w���|�Kr]�k��1v��,"����fP��B_�mM����R��r���ɨWI��T��Vg---�_"E>�K�*{�����i��(7%��`<�{���Ҿ����x�yf�'�O�0���?r�i�:�J��_Gg�C X��-T�ڰ�:/�q���tqk~���a�E�o�˫4�u�~�����d%uV�����z\�sx� ��Pf���SeQʴ>�x��ȣ'qu
��x��iuӣ��u��yt�/Ru;��0Am�[����蝣�(&�|�Ė�zV�'�y3"qwl[������VC��^�.�|�PVy鵵k�"_�~�S�Q���dy!lg~2���A��v]}b޸��D�L��7 Rs����@a�ֈb��Y�)���o�[�o��)C��1��kT�(_o�nn�;J�'u��v<v���Nm���Y���(iDl{U�]9�-ă%	���(48����W~a	���Qתr!��ƌ�8��'��a��/�3g����QC�ݸ�Z���Á��*��<�v�ك�bǢƧ	�͉ւ�V2���f�0^!�V�w ��~�k9��վ��n!K}d��+*��C�p@���L��Y�9b��+� ���)��i9f��rv�.ʔZ�`�3�+�E��l�Jw�^E���R�}�U�)X���:���c���؀3��8�/�`��d��{'�>��b��s�E���˴��V��XB
�͏t�6`fڭ@�M�q~Fz�<���2-V����5;),��K���Z^z��	�sj߱h�Tܝ��P�(����\���$�4x�}F�L�t8����=b*�޿Ֆw�����H��+'''u���à+3++ѥ�-�%��%w�{�'x�V���6<z�r!H={���~���#hgyo03�L-���@��������*�	5_3���:��dL h�O�Ȫ'R"�} g�*(lY5;u��L?m�`z�ժ�N����(<�<�i��XϮ��a��6���^q#�c���,u.E��A����R����;? 	y��sCS��v���k��ʾ��-�Z���9�RNHH���8t�;�G��0�2�^DzBJS��t�k�/��������GX�M�¡Y�ʡ�ȭ�=�E���:����h8���6��>�Z��l~5r(�~@���z(�/��HMi �j���K��̕3�c�w�O�TK�Ǻ�v冗���RPaNmS0��sr6���1��Ws��X����|Z�b��<8c�3B�@�^��M޿Ȥ�R/dG�Ǭ�?9�ә3M��hl�� �or��,���T;���|>�x�"\�\��C!Y�U�l-2����_|{������s'���.��`��*)ͮE�����~;w2xHp�d%!"!{�(�j����DZVا��h��ﶤ�X�-*��������U�a�t#��8�ؤ�ac��A���M��;����?b�P���k��{�2�O�c��J���P�.S�#:�Ԍ�XL���X�^`�]̈���~X�V����M�7=��3QD�Ejǌ�����������Ld�q�C0�D3�ٛ���!I�^薁��9  ��U�2�%pN1�o{~�1�K&�$d��k�m^]�����<Cty�����N������CX^܀!Z����%d�	X�e����4����@��9�S�@��I��7�y岄x�Y�p-��XC�-5ԩ�6r�����zf�3p? CF��G�&�������t�����6 ݳ�a�����/%Le�7����C��D^.�w�9�P����q-a�����+��Y9�\�+�뛱0#6$��M����f�L$� �h�0(��I��g�I� gdU9`���6�3�3�T�}�6�i�z�����YE?j��,���x�I�����N��y 0�	5�K�VaQV�ʠ�(�XRu~Nzhw|���Vlt2�b�J��o:�N�uБlI��s*Ɣ�?_<i�*bn!�2�d"����X�K�m-O>��1PPk��/? W��|�d����ڮ��Y�92)��lڿ{ҿG0��	',5�6{c��vO���\b_�KYf���DN�� ��S�fQ^����oVf<�II$� �T�bK(|��#���sY�¦P[R�Y�*���:f'�Dz�(K��ULx��Eu8ڮ�m�	�l�r���$|.FY�ʪ�n����\_�3��3/�'�V$u�B�M*{@���Y��$`,)����0N�j�
��s;���0�S�`n:Ժ�U�ܮE}�����/~�Y�i�2�d�����I}��V��n�bq�
~�=s�&M���`� �-4�r=]*�</Mb����$�h�uNZ����;9E�]C�&��e�*F�O�]��C脻�Nt�.�Db��D.�S.��Q��k�ǧ�V��,pN0~�N�@����b�I*VBsC��ЕϏ����K� ���Xz��
��dR��L��3M?+�x`�}���׾����C�J�$dΏH`��7.0�!�^Qꤐ|nU�ݲw�L��sC9��Q�;�^�uk�3���:=�/ǝ���Z��m6Έ�|X�-H�7�$��� rg���M/
B7�>�-9;Sw�0û�=�d��HR`�/
�?
�Փ�y�B��{ǆ�R�`�x����=<����fƎ��M���3 ����[4Z���HϟM�y@K\.2q3x����Q����������F��I���EL~��5l=źl����%�I�4ԕ��U`8�z�5w��d�&��S�%Xܳ�Q79}�js�5��h��U�aI�-:y-'����܃D��g�Y�����[�"j�s�|�Gm+��nH5���;D",���9JC���h����Kp���Hm���Ǟ¬��w�mB�����c� ��4[JFrl�e8��͒@�z�r�F�\XR���ӧ��K-$t]�	�P�hiJ�l��u�jz{\)�������q1ۂ�q���c�=�5!t�Е�,���f�ұ�R"�@�"i��_3��氊p��L��Ͻ\] ��t�֧^Z���mP-`����9�a���{l�����v�_�\�~[u7F�`�خ�3�b7�������� %D��;t��xy}�j
.
��Y�.�)$�D��	�s�޳=?��ޓ��M=C�7����F�-���̯)E��)��
�j����R�Y�Z!NE��?j�-�R�����6�� S��ݰ��;1+*83OIV㉹���)�v;g��ˢ� -�`h��al���X���Ě��o~��t�,Rrè����|7B�~^L7�/KV~�YՋY|^�eچ��h�[���`��������^�"���|*��V��l��R�a�W�\�mT[�A����y���ݓ=/��"Mv#�nq[�K�GӴ�Ն/u�������z���J��]ޭW�Z�_��K�6<�M��b�����>�#k�r�y����$8�f�M H%W�dns@?r��D�N�n���R���+#jX��\��� �lv �z���@}������a�X{"Iu_� 1�<0�<�7j�=�5�tr�z���|�6Qh%7,s�Z���?��/�k���c�Y�3de������-�^K<��\��s�-�M1F;P�5�t��h���p0�_�V���������}	ݜ%�R����QG4�\ON�ͷ�<�A�}�lk5ā��{`ƶT1�	�$9|�&dV��(s���	�/#��g�s����I��I|���y��p��+T;�O6.v�g�IۑC_w�8_�p��sM�$��ݻ7���4!����Mv�\;�_"8������f7��d�)��+�����NIJ�孫�e�1�h��"i���T���F��diV2#8;�)WF��x^/����d���%*%�B��}u� �y����>�1����L�1�����%#��r	r2��������}6�_���g�CohyyY��|�.��w�b��Ws�u�kM�3�Ctʆ�EҊ&��'���L�1�i�,q���&��O�	�3����r�PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ��{X��iP  K  /   images/ff54be72-9396-4067-afd9-7c1b32c889e7.pngK��PNG

   IHDR   d   -   X���   	pHYs  0�  0�
�D   tEXtSoftware www.inkscape.org��<  �IDATx��\il\���6���vlǎ�8���',!��&*��@�JCKQ��O[Z�U%ğ��P���DE�P�hÒ&B��4�N�I��3�Y޻=羱�f�č3�`�|�yw��;�{o��?�O G�鉿��T
�,F��I��PY�Àl�r�|*G�T G٠f*+���`�0 T�T�S� G٢a���1ѐZؚ�R$P��"�P�UL�ꨄ�Tq���2K�S5xB�Pc�1��������d&�6
�QTw�3�	��,�dDE1��(b1W�:S����>��ē׉7�T�/4��cě�1�/�|�P,s��I�&����tł���;_�2�G�h��
�x�I�A�-�-��ϖf)f�fŊߐ����.��
	�'�<!�<�'H�Du�����~���j��f}�k+z����U`w�
��^��;K��F�ŝ�0B4 ��¾.���Z4��G?ҖtC����׆��D���i�Y�e�6�/������ð�1T������#G�G�0�Hנ�# ӔԮo�oG��7a�{:�T:�����9��$��M���^�m
{�~���b@�����<0�'�r	������n,�����7�;�ݍ?��"��9:X�R1� Me�.�,�R ����!}!*��^W5zB^�RB`�r���\NQr���&�6��/�'�}�u5\�c^D�t7#��P`zˡ�%4����p̣�'�2t���N���f#2qR_'�ƛol�S�«����;L�䍚(�h��O�1u�T�r��x n�2bK����n2NO�)��2��]']��+���Ε�R��۴2Ϳ-�L����g�h�#�L3n/GU��x[����oa�2|�[����ϛ�ġ�.�G����f�nX<f��,�_�W�=�[����:
�c%��H�e���U��TE�X�p�6���J��*mD�~V�\2is�9���ϨQN�{��YΥ*r~����Y�Te��(����/�C^	��*���+�cPw�SY��/އ�Ʒs|��b/\��1��7��i/������s蚂�ZD}MttP�[p�#>��b�1n��iS��Q":gN1����l<FLT�j(*�ʃ����6d�����R9��I�zq�m5x�߇�5�`(+	H���?h���܃=WH�SR"K�wei@2{ Ew��������4��� �z�r��X�\�7��P��0�yI��O��`��q�K�k��5�m�q�kv�<��y~7ml���-m�#��,�p�����C���Ç"q,_R���81��儬��]W"5�rv�$�Զ��#R�>w.�)Ǳd���@`���y�ĸw6Ǒ�N���;�"�i�j�a��*�plk��{Z�|N9VR���M��ה��d!���i�o�l[�5�#w��3q��P|��S|���j��q=fNϧy�q�
+V�����w�p6%�:3:
�*��2�\:0x���{��T���b|��7no��7J��(�ó�j%�_x}���������5���kh����^��Ϟ�%�K0��.�b෯���kPR��/_�T2��u˨P5ݏ��y���_?s�y'��:�޿ �y�Uy�,<��:y�x\H�[{���B<z�<� �Z���5���)~<r�\<��6EmA�uI�V����?}�F���;N�3o���kN�@[� ��L���������@�l��%�Ȕ 
)��gL��<�����:p5������+���#g���)m]�CXD>b��)���b�Ԧ�E`������jƬ��6�؟���PT�o!�h�$3�v_ɇ�uؤ����y�/ _9%@��'�g�`�_`�+��m�m�h~c�4n	ǂ+�IA	�f��ɹ�'������4�l	&#>Ի,��;�U��`�������#+�N�aӮ��bS�rY1�;?o��p������X�7F ��i���s��;�Y�!��,�a�t�!�6v�d�?^{����v�[ 	��m�l%�G����	��\+��mn�>�l��a�	t������X�t���Zۃ��Y+%%8,�z����K����&d2��I��dY�Q�r��#ܾ����M�>d0��Zq����F�������
�USf��PU^ �v��Vɤۮ��~�$�@>0;K6Q'[���T��+����hEiQ@FzX�I�(��Qo���7�������E�����?Տy�S0��X����
S$���F�?�&�d������X!�VO`��FuyiR�<#�)���C~� ��}���c2 P/�	e{���[���H��B;oH���Jں�d4�S�H<ž#�h8�Ѓ��ݲ�c��e�鑼C��l������Q�x������Kec+�h�R6�9�&�Y��퐟9l1�O�qlj>�3����#s�>�&�ە�#J�f��&{�j�;�5������;�G6�{��zEu�T�����L�'2ַöQ�Re~b�T�R�i�pD�v��4�2�0e>!%M�y��X��8�?��LeI���
�/�F���1�t���s��˴} }J�*ι8*��T�g�?(:_�8 9����2� ��D�r���I�(V����
{6�ux�8�3d�o�y��1�e
ѴH?�w�CKd�|-�Ɣ>�Χ���G�J��s9�\���q�1u��2�Zv�g�I7SL�2N�<�};�b??��g�9�d<I�'O�����sL|>�_P��0ׅ�)M���=# %hZ��6�3���/�D$����SNӻ����my�4b�]tůfN��o&���P�%�����i�g����х���-MF@"�H�E�M��K~�7m{�@�Ӟ���|��CCCC���ԷN������P��U����N�1��I�E����n�1��þ��<&^#她Q@(11]~�-}�w�HA����^T�R�0�%E�4Û���3�C��k�����dc�]5��FKsy�/���ϓ��V`��� qß���`nN����?�%!/��W���DZ�d<���>*%p��'Z,�C��=&�]!�qw���P.���<A#��w�G=Jr��F}��o��xBؙ����1/:8s���:Ge�԰(T�gpyЊD�� j�?�Q	�E�	�[=�|1�*w$*�a�r���q�V*�PY29i|D�.1��烰�y�������r��e��"�f0��bv���KAK����r��``Y    IEND�B`�PK   +��X ��ٚ  �i     jsons/user_defined.json��n�F�_E��.VC̜��?'N[c'��t�"(�+��.��Ah_f�i%9���(�E����(�7C�|�2Q��ˏi�h�Z���1�i��x2�5�Ӫ�hA�k+_o�?���՛Sw^�����h�)�#���x�;�L��G�a�b��X-��&�v���<Z�Wi2�⫱u^
2�V(� E¹�D3�������{q�����r����/��K��".�$�iG|�X��c��`RqQ�����*7;�,�O��VA�&.GKt`�C0�&}�ӹ{��Ux���g�r�sp�C�O/��I���O�ru~<]\���'��ܘ�BXE)nv�٫�����it#�9ϫr��
��<�g��[�RoP-�u�ϧ3\#l�@O���� �����9�|u�gΧz��'�Ɵ'��[ݮ�-�����7叏:�[�э>�{��>yҩ�w�Z_��ٹ��������Ux���r:Gs�����E�/�kp�P�_Te*�o�xau�n�q��k�F?�αW��ȕq�:���[��it��E5��I���|T*h� -;�$HO	H�w�ra��͐#�눼�L���0�9������OYH%��Ҕ8e-�;��#��y���V\����fW�&�~%}����������1���sp�o�u�DF��C#sv����nU�Ϊ�l���.�QYo�We��m7�h��e��h�H�H��(&����t&�����.�� �
�˶m�m�((������J�&�vwV
�ǸwxӖ` ��m��}l��q��8;���6�0�3��h���)�Pl@��m�+N�l^c�
vX�܃�OW��b�<�����
�l����)a\�}^n!�P]�(� �_گy|;]L�,}Y7O��֍��>�6]��.���o6������Mb�d!G�b� ����f����j�u�����N��UB��8���%����,(C�疤��0�*a�bY�W}���ĴW�Й%N�B��L�,���j�~l�ue�>���se�3�ZJ���W�~&):�*0�q�d�Sc�D0^.�A�m����/�� y�	��`����+��I�h�����u���ժ��I��Z�:q��V��9���@���L���&Ljw�1'ۗ�w�7]d�ye���W��}���Ń&0?"������^���\%�� eMb ��3Fg�P����Aҽ�F��|�
�z���O��ZAr�!I�z�*@�`�P�ykF�y�l\����	�	��B����J`��I]0�]$oɗ��^{���7���^a(VK�K0�%̯����u9��.Ç�k����3<�.�W�݆蝴Q�H�՚�c���R��b�L�����IzOL����hH��NX��@w���]J�%�*~����︪��)�_����4#��7��6"<\Z�|���ʖG'e\��`�87Y:�%j7*"��5�1��z�E0�ﳧǏF�/�^��_?�٬����6Q�e .1Z+��S�9�D�d��:BHŢ�i"��C̄�:91ÊuVI
Xh�&�{)\,�|��%Catm��V��رv�����C�Nb[�°!K�t�z����Aϕ�μ��Dڂ�cim�M(�ֻmy=�~u�ߓ��=����[p�x^���<4��4d�:	I V'CMp��c�H<�����]���f�g�)A��1�	��<�X'z���F&!�ǟ�'Y戵"�rA��AY�T��X5$��J�aZ�q�z�+�K);��գy\M�j����x=��y��ZΫ٬e��fZ<z)(��a-(��bae<�5Zj!�oZ�DC1��A[�U�#�&Z'U'���:�_|��6����:�*�}��]�d�fv��4����n|ߜ�9{z��&�e�px�����#��d_�EZ2,�z��=h4�����l1�4w�=����jQݬ�i/ѷ;*"��^�G�S�65;��ɺͿm ��(t��s���#�-�D
�����m�L�Hv�6y��N`l�9��(�Sv����'{���&V��5��oL��=f;���}e�A���%��vC-AK����/��tOYۭ��LOUӭ�dl����n�&c�]�^��[���:�Q��2��xO�n�-�K�T��ZB���Mo�]��j7\�%x鞪�k������JX`KA���Xo�����h�X|_��(ʎ�bR�o2�)�"{��
3��b٘���-�B����k$��w�*�&R:I�YL��o��w"XJ���g8�K,PnU6	��Ҷ�r_9�Qώ�2��=�@@�l��~¾�H;�>zueO�ޖ���>��>#�юX��Ͽ���~\���9:�/�����1��y�m��=��+���?�I=�D�ݠ+bgbuY^7���v�c�|S�-�����^E��o�n��?���/���@��z�7��s��y�ؕqq�'y�Cb"'�W[��[x���Dh��aDn��8�%��5xc��G<���0x��#a��G<���0x��#�~S��K{'X����z�\;|�L&9�dX
�7b�9��Z T�Ā2D�舋ɐh#�!�l&X�A'Xi�M���{M�r�q�r&L%U�M��%��S��4��!v�{��C���c�ǣ���2�1O�K��8g41�r�����۹(���sB�ç������Y���-߈��!x=֒��������cԁ�@���G(|ʄg�`!R���������������������������������r�~�F�W����N���k:�-P1"@Ib�bD�艋`�1(���A�3���u6x���d�I
)/-���)V�ط,����4�TVs
�ßWEi���0���E�&�G�g]u��Z^�{<v��?9�0�$���<�&��4V3"���$2��X���>�PK
   +��Xv_��9  	                  cirkitFile.jsonPK
   ��Xyɜ��  �  /             �9  images/110f4c69-ce42-4daf-8800-65b9db14e3fe.pngPK
   ��{XR�/�+ �/ /             �V  images/12438572-56ec-4fe3-962c-a8f31caef061.pngPK
   ��X�䓶� � /             ɂ images/132fbcdf-34e4-44dc-827d-09a965026955.pngPK
   ��{X A��?5 �J /             �6 images/1a82a878-f7f8-4e20-9f5b-ecefcb5937dc.pngPK
   ��{XF&�!    /             Xl images/24a54a69-5cbe-4d66-9ad9-6bf107554def.pngPK
   ���X��g� 
  �	  /             �� images/4f5a6b59-a216-44d1-a198-112719b334c8.pngPK
   ��{X����?  [G  /             � images/55b8074f-3515-417a-bf4d-91f9a1b9fc8e.pngPK
   ���X�?HU!  B#  /             � images/585092fd-6de4-462f-8499-92296fb2c536.pngPK
   ��{X�c^��  �  /             �� images/817a53b6-1ac7-4961-8971-5b4538e0cf16.pngPK
   ��Xd��  �   /             � images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   ��X�1.:�  )  /             �4 images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   ���X�� �f  y�  /             �S images/96fabd4d-0b16-452b-94e2-688cfcbce531.pngPK
   ��X?S��� 2� /             � images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   ���X���5�  1�  /             ��	 images/a437e5bb-8d3f-4b3f-8093-72e2f97ca498.pngPK
   ��X	��#u } /             �'
 images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ��X$�8�l  �  /             3� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   ��X+L$��� �� /             � images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
   ��X����<  �  /             � images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
   ��{Xw�'<�  �  /             �� images/bef45656-42b5-4670-a699-453aaa19c38e.pngPK
   ���X��g)�
  �
  /             s� images/c1fb8ae3-abb7-4800-a199-c8a1e0562abd.pngPK
   ���X$7h�!  �!  /             �� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ���XXs�銙 � /             �� images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngPK
   ��X�GDU7� �� /             �� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ��{X`�/��1  �P  /             As images/e80f2fa1-d37d-41df-8a09-120fd0c34151.pngPK
   ���XP��/�  ǽ  /             #� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ��{X��iP  K  /             uW images/ff54be72-9396-4067-afd9-7c1b32c889e7.pngPK
   +��X ��ٚ  �i               e jsons/user_defined.jsonPK      �	  �p   